�� sr gui.PlayScreenK��0� L 	inventoryt Ljavax/swing/JPanel;[ inventoryPicst [Ljavax/swing/JLabel;L m1t 
Lmaps/Map;L p1t Lmobs/Player;xr javax.swing.JPanel]D
��B$  xr javax.swing.JComponent3�c&l�� F 
alignmentXF 
alignmentYZ autoscrollsI flagsZ isAlignmentXSetZ isAlignmentYSetZ verifyInputWhenFocusTargetL 	actionMapt Ljavax/swing/ActionMap;L ancestorInputMapt Ljavax/swing/InputMap;L bordert Ljavax/swing/border/Border;L focusInputMapq ~ L inputVerifiert Ljavax/swing/InputVerifier;L listenerListt %Ljavax/swing/event/EventListenerList;L 	popupMenut Ljavax/swing/JPopupMenu;L vetoableChangeSupportt "Ljava/beans/VetoableChangeSupport;L windowInputMapt Ljavax/swing/ComponentInputMap;xr java.awt.Container@�s�' I containerSerializedDataVersionZ focusCycleRootZ focusTraversalPolicyProviderI ncomponents[ 	componentt [Ljava/awt/Component;L 
dispatchert  Ljava/awt/LightweightDispatcher;L 	layoutMgrt Ljava/awt/LayoutManager;L maxSizet Ljava/awt/Dimension;xr java.awt.Component��Y�<�� $Z autoFocusTransferOnDisposalI boundsOpI componentSerializedDataVersionZ enabledJ 	eventMaskZ focusTraversalKeysEnabledZ 	focusableI heightZ ignoreRepaintI isFocusTraversableOverriddenZ isPackedZ 
maxSizeSetZ 
minSizeSetZ nameExplicitlySetZ newEventsOnlyZ prefSizeSetZ validZ visibleI widthI xI yL accessibleContextt 'Ljavax/accessibility/AccessibleContext;L 
backgroundt Ljava/awt/Color;L changeSupportt "Ljava/beans/PropertyChangeSupport;L cursort Ljava/awt/Cursor;L 
dropTargett Ljava/awt/dnd/DropTarget;[ focusTraversalKeyst [Ljava/util/Set;L fontt Ljava/awt/Font;L 
foregroundq ~ L localet Ljava/util/Locale;L maxSizeq ~ L minSizeq ~ L namet Ljava/lang/String;L peerFontq ~ L popupst Ljava/util/Vector;L prefSizeq ~ xp               �           R       psr java.awt.Color���3u F falphaI valueL cst Ljava/awt/color/ColorSpace;[ 	frgbvaluet [F[ fvalueq ~ "xp    ����pppppppsr javax.swing.plaf.FontUIResourceBć�"�G  xr java.awt.Fontš5���Vs I fontSerializedDataVersionF 	pointSizeI sizeI styleL fRequestedAttributest Ljava/util/Hashtable;L nameq ~ xp   A@         pt Dialogxsr  javax.swing.plaf.ColorUIResourcekS�����  xq ~      �333pppsr java.util.Locale~�`�0�� I hashcodeL countryq ~ L 
extensionsq ~ L languageq ~ L scriptq ~ L variantq ~ xp����t USt  t enq ~ .q ~ .xpppq ~ 'pppsr java.awt.ComponentOrientation��E��c� I orientationxp   ppx        ur [Ljava.awt.Component;��u  xp   sq ~                x          R      Spsq ~      �@@@pppppppq ~ 'q ~ *q ~ ,pppq ~ 'psr java.awt.DimensionA��׬_D I heightI widthxp   x  �pq ~ 1ppx         uq ~ 2    psr java.awt.GridLayout�#��K�� I colsI hgapI rowsI vgapxp   
         pppx           @	  pppppsr #javax.swing.event.EventListenerList�6�}���D  xppxpppw    xxpsr java.awt.BorderLayout�ב_ps� I hgapI vgapL centert Ljava/awt/Component;L eastq ~ >L 	firstItemq ~ >L 	firstLineq ~ >L lastItemq ~ >L lastLineq ~ >L northq ~ >L southq ~ >L westq ~ >xp        pppppppq ~ 4ppppx           @	  pppppsq ~ ;pxpppw    xxq ~ 4ur [Ljavax.swing.JLabel;��%i*  xp   
ppppppppppsr maps.Grasslandsw��|cL�� L randt Ljava/util/Random;xr maps.Map9��M��� [ gridt [[Lmaps/Tile;xpur [[Lmaps.Tile;�g�ߢ�
�  xp   ur [Lmaps.Tile;}�ߌo�>�  xp   <sr 	maps.Tileu�%q�mx I heightZ walkableI widthL itemt Litems/Item;L mobt 
Lmobs/Mob;xp        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psr mobs.Mob�����C 	I armorI attackI 	directionI goldI healthI locxI locyI 	maxHealthI speedxp               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L         psq ~�               
   !           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ͉PNG

   IHDR           szz�   �IDATx�c`h�  ��ve<㒣��r���2d9�9d	[�*�-�}o0#E�f ��� �#i� b��� �,dh� p|�j�#hf!rb�i�G����4z\���8E�D��.z�B�~tK���G�(�`��Q0
F4  �+�'	ŧ\    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw�   ɉPNG

   IHDR           szz�   �IDATx�c`l`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R��	X�4�`d�	l�-M�B	�n�V��AbV�9�� ��71e ���2�f�=
F�(�`��Q�  b#����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   2           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   2           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw�   ɉPNG

   IHDR           szz�   �IDATx�c`l`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R��	X�4�`d�	l�-M�B	�n�V��AbV�9�� ��71e ���2�f�=
F�(�`��Q�  b#����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   6           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`L`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R�8L��r a��� �S�D9�-G��h�͖�`��Q0
F�(� ��$8I�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`L`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R�8L��r a��� �S�D9�-G��h�͖�`��Q0
F�(� ��$8I�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppz     {�PNG

   IHDR   P   `   �k�   BIDATx��=��D�{/!��D@BH2/"CD$oH���F`1,��
�p��9����yvۖJ���������v��k��k��k���m�|�t�q����_���v���o���5��`5p��k�ۈ}���H����7�Á ���� ��F����k�y�p1�f� ��s�F(P9�?,H�wJ]K��yhڬҸQ��CAx��m4 `X�
:G�C�.*f��I��.��Ѵ�B4-t���c�8���@0@U\ ��n���f��r>������5����r��x^՜�Q�P"C�.���"*�kY��q��
��-��p`�MrҚ%��ڙ�Du�M#3�G�&��l�%>V��7�l�KR����}#
��|�Ξ1T�R�Q���S���{�\��}����p��� άD�k���t��˾;*kU7bn�qlҕ�e��f(O@T~L�IV�w(����"�L[��`p��Kw֔})Ȭ	ʍ�-R��	fQ1*ʮI��}��4eQ��5~�:�����T��k�T�p�gr����R^Qb�Z���R���hB�JrU��=��f= ���FT}G��f5�ڑ��9��y&G� 1e���^Ư�1b��Y�:W*`�]R��&:K}��\�r��g*��M=�S��̵b�KL]AT�W3 *K�@E�κ��bթ�&��"�ʸ�2ۄ]�KBl��A.�����L�&��sTٯ����z� {f�,���6,TMms� �={RIj���2q�N�P�TS�P�X�/t{��P+v3���y��J�^���%�za" ^�S-���U��jy��y	 ����>ǻ�%8Х2K|�� �q�� ��R����r�έu`�8�	wK��6��}"�R@�ܳE��dF�+�;y�=�X�m�w/Z�䨌usf����ΪKY��+7C�����Em~�L�+�Z����rOU�T�z  ��n��D�J�*�-w�\���V f%!���u��"x���E���0�oԤ��~����؄���~(�9�%�;�B��kz+lY�����JIן���)�25�T�?w�Q�]%�SՏJ�\��|?p4��s<T�Q���9�Ytu�|6����f�S�P&]�jؔP5�ϔ�Kq�z9�����3(
�:�%��=����]�w���_��&O���B��5VL�݌^y�L3��&�˒�
�j2�f�&�)؁W�2��)�H��7�}��}��%�8�����Y���"���W���yf�c�Os7Ae��o\�������?~�d{uf�S��Ο��\�{�0������k@\�3�;��+f�0���s�ʻE{��*���~Ϫ������?�ŵ<7v�?�1�P`��"�M�^�����s6-�^b� "\(�����Fd���#�?5n�:ש��[��!*�����x8p���`�:N��#o1I�C�h���ۙ6��Pq#,�2��vƍ!*�f�PN��ۧ�rP	��`qzx/ >i���y�#r��!�`��Е}��>=�o�\Gu�*�f����z 1T�����l�T���_�� T
D_x����;VT�@.��w��KѴ;�ćU������D vq�c�0�����V-+�*Su��W(���`T��q�� �҇���	�ȩ@;�a�ǭ/չ�yH�m3x��S-}u.��S��A*?ŵ���@����8��c�����멊!�5U�ͦ�{su��1�z'�j��-wd۲�G%y D�ɠN��r�a��̒sܺ�h4e�>t�����۵��f�^�A���um��b{�ҥ�<|m    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`L`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R�8L��r a��� �S�D9�-G��h�͖�`��Q0
F�(� ��$8I�    IEND�B`�xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   1           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ɉPNG

   IHDR           szz�   �IDATx�c`l`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R��	X�4�`d�	l�-M�B	�n�V��AbV�9�� ��71e ���2�f�=
F�(�`��Q�  b#����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ͉PNG

   IHDR           szz�   �IDATx�c`h�  ��ve<㒣��r���2d9�9d	[�*�-�}o0#E�f ��� �#i� b��� �,dh� p|�j�#hf!rb�i�G����4z\���8E�D��.z�B�~tK���G�(�`��Q0
F4  �+�'	ŧ\    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��SK
�@-^E
�����Ap��#x��C�"�=E��yC��*�ȃ@H�L�-	�vԿ����a��$z�~�ו�t5 �M�`ξy
 !R`Bh�3qI$d_"
�<�*b�?�㶚ׁB�Y�-�݂�aI3�$�~�$V ��W��c�)X�n�V�������m ��N���W`_��N$�D"�X
^�45aO��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
               z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   0           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L         psq ~�               
   1           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ׉PNG

   IHDR           szz�   �IDATx�c`l`���dLw���,C�ts�"�����w3���d	� 6H�掀�d!�ݦ� 6H��!�%�t�RCS����i�0-U���0z�YN��	K���=a�B[��&Ll	����0A&O�f1]JF\	����Q0
F�(�`�z �/7V�@�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppwW   S�PNG

   IHDR           szz�   IDATx���   � ��nH@   �  ɵñ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   9           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ɉPNG

   IHDR           szz�   �IDATx�c`l`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R��	X�4�`d�	l�-M�B	�n�V��AbV�9�� ��71e ���2�f�=
F�(�`��Q�  b#����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   �IDATx�c`8�|m��Ș��Y�����E����f�7��Al���9�B0�M�Al��C�K�%��9���@t�������A=�0L�n	f1] �� Y�t��(�`��Q0
F�( �G�M�~ʗ    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   rIDATx�c`���a����t�d���06��v��l9� ˁAv̓�RU�?�1莢K� 9�C@���r�(�YN� r �,����|��Q0
F�(�`��� @;ost��Z    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`L`���tLW�R�?�x
��l<���! �a���m8F��#� �5�@|�;�RU�?Â�R�8L��r a��� �S�D9�-G��h�͖�`��Q0
F�(� ��$8I�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  
  �PNG

   IHDR           szz�   �IDATx��T�	A<lE?~�s5X�`�`b-��*"�0�{��䕁p�l&3s;�����!���J'�o�q�Za}8�$�¥rݵ�$�DۋV�`S|��/�\,`c==��[S($�(L������Y�Sz���ލ��p���Pg�2�,�
��߂�Iј
��6X�ϲ��>��1|��p�`��B�U(
�B���o��bb|    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`,`���&U�,������9
��@|��T�8 d�0C���8����L�� �A�RU�?�w �&Y�1��ɡ�U��w`v��� 1��0uTw ��� �4s z(`�=9��( K�	9!"�iZ.��l����(4`�W�[I�+q���'� �FO�Ri!'��9�'�(�`��Q0
F�  �,EB*ރ    IEND�B`�xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��T�	�@<lE!��`� ؂%؆5���� �ӧ��d&���=�c�\v!;;ٽ�~Ĺ�f0���c��Gk1�����+@;R�<�� �e��u�o��g�(�u�#v���|Z⌘:�d���� ��/�	�.�{<�qb���C����迆�^��t�f�ښ�a��Y�_-3�6�V�w`/$7j�-��څ��
��(�����
~�u�+8�@���=�O�K_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��׶����4w��$��0�����,F�[�*�-�9 ����4��@v HƦy(�,Y
�.�� ���#Y��KN�;
t��b�(�`��Q0
F�(� /��(    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   9           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppz  (  $�PNG

   IHDR           szz�   �IDATx��TA
1,~Ea/^�7��/���o���"=
ޣS	���x��@�B3I�-��i؉e�F�R&���x͕��\cw!�T'gRP��z�M�<O�B- Uk����5;c��37X������ b��y�g2�r�W�3Y��k	༑�ް&u�5�}�.�v+�v5^��r$���k�tB�U2�@q!F���>T ߸5 ���pl�_�F��D"�H$�/>�4��!�q�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   �PNG

   IHDR           szz�   �IDATx�c`j`������6pLW��-��`���9 �OU�~<�����Y��w3Q��`˿l<���� ��b�#� Ñ-G�K �qtw r��
4��6��Mr���>F��@�Fv �OsX�*�aXp�[
���K�Gv�lJs �)r�d�`��Q0
F�(N  	�&s ���    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx��1
�PD?�F!MZ�����B�"v�/!be�	��ERXd�b���|x������:W����n���bϽ5���{��Hd>�8�0��h��`��H�ˍѱj@������Ə�է� ���|� ����;@�,�4x�Y]���^�A�M6�؍�� �������)�(�Y��*%��+-�T*�J�R)��G@1�����    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   |IDATx�c`X�|m����m�ħ�����0�a�ǧK��Y��w3��y��[`�
���� Y � ���$��� �Z�,U���9H�n� �0LW�G�(�`��Q0
F�(�7  P��-u�g�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   xIDATx�c`��  �?���pG����H`�8�#[n��L߃,���:@�2��n��BX4��4O���GN|�耦�: d,�aQ ��މ9�$��Q0
F�(�`�  \���᧵    IEND�B`�xsq ~ L        ppz    �PNG

   IHDR           szz�   �IDATx�c`x�|m�� < ���Ï���.�Y��������׶�; ����!���`K�1�b��`�a�:�9 9�a�<���x 9�pL3�0< � ��-���_�q���x�:�3��งaP � ��,�a�9d�P�% �� �CzX(Q-*�-Gw�rZ�=�Q|u ��4s���H�D	�qTzbCf�h�8
F�(�`��a �8I�#��    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
              z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ��PNG

   IHDR           szz�   uIDATx�c`� ��m���b����?��/O��4w�p�� �_����i�d�|�� ���TU�°�F�$SC󴀜@ħk.��9Q���`��Q0
F�(�`� 7����jE    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   PNG

   IHDR           szz�   �IDATx�c`8�|m�� ��Ms�M���������bt񽥪2�B��1M�M�d��al��9��Al�YNL�#[
��s�XNJ���rG@�
4�st��s����9VG@C����;b@,�`��Q0
F�(�  R{���_    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L         psq ~�               
   )           z  o  k�PNG

   IHDR           szz�  2IDATxڭW1�1M6�{�~����˿SP=�섯"|�"�؉
�6�o-�~!XZ�X[(ba!ZY���haa)،;�3�\.��ăw�f'���IfV�"h�W���A٠h�50�_j���T����JE&��g%:���ݤ(��,2G�4�9�	脅�XH�׉D|VžQ��J0'�MqQ,�\���d�<�����C�?_��j�oУ�����L߳�9=�NJ`/�3���10����D��U�.�=�������$����3}�[�Zȴ�6@eO���ow�gZ�r�ߺF�Y�&�V��T>^=
�nٖǬ%�c��?ǌ�ŀ�-Q&�J�?~�~�-� WLRO�J�F�"T�;ŝ�ڰ���� �d�2v�."��Ң�P�� >�܉�	�;!���ʚ�}�V��8?�ZY� �B�0
T*��؉� ��7�;J%§,��Lwj�&0�L���y�R���Ĳa4	�BlV�(�[ivV>82��.��_/�rF0i�0�<D¶�_�}�U�$�h�tA,}�����*����Ö�T].б{`��3��g"3VP	 (��5A��3qeZ���=�u	��ux��~T,du�(�/+!��jΎ��`�-����s-��+X��@Iw?�r�`���$|v�(�r_9��^�B9�7�"$s��"��^̝:��}"�* �2���Dg���h#Z�JHVLr�hSJ���X;1`ȗ#�5���%��L�ߴ!�c)\:��;*ܔ��m��sO!�/����Jr�qI���E���W"EW22���A�x�|оZ �o>�ł������_1�n��w    IEND�B`�xw�   ЉPNG

   IHDR           szz�   �IDATx�c`��k����m� >= �"t�����0����rt��Y��w3��y��[`�
���� Y � �all�"��%��@�Z�*��k�G�Z>��<��+�h���/Ҽ �plqN��O�0LW�G�(�`��Q0
  B�W�&z}    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw�   ݉PNG

   IHDR           szz�   �IDATx�c`��  �?�������=.��#@��Y�D�,U������ā����Ā��`�
�F,�0<J�+@�,DN��(�y��Ys�ve<�RX����4�}	� r��h� ��Fr�����Q@�����#�j�(�`��Q0
F�� �ɥ���w�    IEND�B`�xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xuq ~ J   <sq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xsq ~ L        ppw    xz     ���PNG

   IHDR  �  �   [���  � IDATx��ݱ�%�-�t�k���8@�*�h�7a �C(3�@��7�yW;�4�U���Zv�����?��������?��������_���������_�����z4_��~f���\��ܙ]�<<<<<<<<<<<<<<<<<<<<<���e�{.�Q�����l�E�QX(y�e}�����=��ki7������A��ެ�,�3<'��X�eK�A��|���Y�I�Ѿ��yxxxxxxxxxxxxxxxxxxxx>�s�	�x�����������D2����w#|�z!�3<g��tw���ed�������o�gxN���3��w-�e�7�ѳߓн��������������������������n�����x'��:u��e��N�<Oc�}�x�*���lU�vw�;ĺǰ���r�Ż,�gxN��h����;�}x�6ݧ"���!6�����������������������4��N��Ǿ����cU�;�wg]����&��zΊ��+����׾���;��/2�<<<<<<<<<<<<<<<<<<<<<�����MY��Y=�I ����_��gx�����r��Z?տ~�w�Ѭ�i�g�Y؃�V���D�O��)����5V}G{���i�)r���^�)���������������������|��t|EPg����޹!Y;��ۑY������������������������t�i��P��էe�M�����w���w�gx�j���Q}�[������ai����������������������<�sz�z��5w���z   ~�����6���J���������������������y��?�a�du���3ȝ�yZ�w����~yv���������������������y��|�]g��+�z�O;�o�g�{}U��8f�gxΚ�^Q ��4���s�����5��'-�{��������������������������J�﫧��ջ��`����GҒ���������������������y��c�����w�W�Uj�t�H����������������������� �yw�a�E�M�2��Z>������������������������h�y���L�;	֫zG���u��y>�sI�cxxxxxxxxxxxxxxxxxxxxx>�sR(E3��I��qW_a��k_�u�)��\7�3<'���x~���i��1��.�n�������������������������7��a�a��B?�c��h^k������������������������I:3�+O��v/������g���k�gxN�_f�Ý����<�<��f(IY����ܙG�����������������������t�Iў�����'}Tw���B�f9]���wd-�3<'g v6G�$Fz.r����>������yxxxxxxxxxxxxxxxxxxxx��9=b�m�4�;1�g�S��S6��o�yxxxxxxxxxxxxxxxxxxxx��9����d;�Y�z�������w�'�?Z���������������������<�s��y�6Y�.�ˈ�ަ7�F{:�/��8�3<�׬�{{���Z�3}�^{�Ꮑ�<<<<<<<<<<<<<<<<<<<<<������t_g�zE��y��2�v{�L������������������������y���ޝ�Fx��t_G��$���a���F;�G{δz   �3\���>��N��	�n���wr�.к������������������������s��8�0��I�N�t���8� �����@k�gx�T�I���t�̣SqC��������������������������y��w�g���)�����|�ܿS�W���x�gx~7�� v�[w��Ч�Д��v'LgI���}<ϧ{�h����2lq��_�R��4�{�:~q�*2����������������������<�sVDt4Y���%=$��=�|^�B����"�8E�x~7�������N����T�zJw��í���_���n����������������������<�sҺ����Q�?��;ˣc>���F\OC�}�"�G{Nؙ��5P��8\��Q����� ����������������������<�s�	�e+ѣ��Y����4�S��������<<<<<<<<<<<<<<<<<<<<<�9�<}��g�w-�F������	�.������������������������8��MK�Ar��Ȥ��h_��<<<<<<<<<<<<<<<<<<<<<�9߄}�li���cҩ�w�dH{���F���B�gx�,^���j�-�/��z9���}�w��<<<<<<<<<<<<<<<<<<<<<��Wwg���Z���o>�g�'1$�{!�3<'	�_��9�N�u�dy�2��6y�Ɣ�<<<<<<<<<<<<<<<<<<<<<�U��9z٪�-��w�u�aOٙ型wY$<<<<<<<<<<<<<<<<<<<<<��\u�Lk/qw����;m�OE��/�Cl4�3<�h@ߝ�5�}W���Ǫ>w��κ���M�����EWp�]=�}�w�3�z   +^d�yxxxxxxxxxxxxxxxxxxxx��9��q7������z�� 2��B�0?<<<<<<<<<<<<<<<<<<<<<��;$��{���~��^�̣Y�\����;��噉<<<<<<<<<<<<<<<<<<<<<��9+R:�#Ϋk��������S�~m��S����������������������h��������[�sC�v:�#��z�����������������������Ӧ��/�O������M��L��;�<<<<<<<<<<<<<<<<<<<<<��������
�Ή��S���z���������������������y�����:1k��?���]��kme��6�����������������������&�����.qW�f�;�����9T1������������������������� �����4��W�T�v��T����>uq��.<<<<<<<<<<<<<<<<<<<<<��5M��@��i����U���kx�OZ�7� 7�<���*�WO���w+=�"�s珤%���������������������� �Y� �#�U���絛j���� �ޅ������������������������L�&���+�zeZ�|�z����������������������ў�~W��w�W�����:��|F������������������������|��P�fH��>:�㮾ª�׾��S�n�gxN�1\�����! �&�c��]��\7�3<�o&�������~t�Z�Ѽ��;%�������������������������tf�W����^��i����x7�=�<<<<<<<<<<<<<<<<<<<<<��T���H�;-�y3�y:y"��P�0�b�睹3��l����������������������鞓�=)ݽ�;O���X둅��r�b7����Z�gxN�@�l�4�#H��\�:EW}k=�z   ?Z���������������������<�szĺ��i`wbt�Z���#_g)�l���Z���������������������<�s����v�;�>�lӣ��;=�|O:�����������������������y����	�m� ]�!�Mo֍�t�_Zwq�gxN�Yo��:*1%���cg�:��|��yxxxxxxxxxxxxxxxxxxxx���G:m�Δ����?:d$����0�5�������������������������;$���龎��I\�~hݍv����iKg�:��}|�27Vݠ5�=���]�u9�<�>!q.:a:��6����q�Ad��7��<<<<<<<<<<<<<<<<<<<<<��ؓ�m��T�G+�:�����/h������������������������t�fw/<R"�'�������\���"<<<<<<<<<<<<<<<<<<<<<���n@����h��O';�)���N�Β<],��x�O���$�ce��dK����i���u���'Ud^���������������������y�笈�h����JzH6�{���d�t��E�q�<<<<<<<<<<<<<<<<<<<<<��n@w3;�͟�N=M�8���nw�[��׿ ���t���������������������y��u=E;$��s:�w�G�|tg}������E����4�3w=k:�zq�B=֣n��-�5~/���������������������y��$:�V�G�ų2ﯧix�H?Z	#�͗�yxxxxxxxxxxxxxxxxxxxx>�s:y�ni�~�Zڍ�3��}���]������������������������q�-���v�:.�ǑI�Ѿ��yxxxxxxxxxxxxxxxxxxxx>�s�	�x�����ǤS��ɐ�j�ߍ���<<<<<<z   <<<<<<<<<<<<<<<��Y�:��վ[�_���r��7����f�yxxxxxxxxxxxxxxxxxxxx��9���tsߵ����|F�~ObH@�B�gxN:���s������eN;m�<�)�yxxxxxxxxxxxxxxxxxxxx�9�h�s��U�[����Þ�3�=�Hxxxxxxxxxxxxxxxxxxxxx��9�ꢙ�^����w�t��ؿ_���h�gx�р�;�k����׏U}�,ߝu}�/�<<<<<<<<<<<<<<<<<<<<<��9+:�����z^��kW�g�W��x���������������������<�s&��nT7e�O�e�'d6Z��~a~xxxxxxxxxxxxxxxxxxxxx��9w H:���y�k�T���ޙG�6���-fa~wX��3yxxxxxxxxxxxxxxxxxxxx>�sV�t�G�W�X��qW_�%�����z�����������������������ў�-�A�����z�d�t�oGf�;������������������������=�M/C=^V���7����>ߙ�{w�yxxxxxxxxxxxxxxxxxxxx��9�)~s�E�n�ק������������������������������u0b�������z���<�v+m������������������������L@�Փ�]��� w�i��	�s�b��ٝ�����������������������uw�i�ۯ�>�𿩞��U}����]xxxxxxxxxxxxxxxxxxxxx��9k�zE�7��/��q��z7���v���o�An�xN7�(U���&wW�Vz�E���IK�������������������������AlG��z���U_�V���"��<�ݙ�M��W4�ʴ�k��;�����������������������=�e#��2��$X�����uz����%����������������z   �������t�I�͐v'}t��]}�U��}9�=�(�s�<<<<<<<<<<<<<<<<<<<<<��c�Z���?�C@�M��X����n�gx��LP��݇!��莵Σy��wJ�3<'���H�<�۽4��n{ߟ�n�{�yxxxxxxxxxxxxxxxxxxxx��9�~���wZ��f��t�D֛�$ad�Z�;sg�ق����������������������='E{R�{�w��=Pݱ�#1��t�n��ߑ�<<<<<<<<<<<<<<<<<<<<<�𜜁��i�G���u��&� :�z�����������������������y���u������螵N��G��RL��׿	����������������������y����1�$wd}:�٦G��wz���t��h���������������������� ���1�dA��/#Bz�ެ�頿���<<<<<<<<<<<<<<<<<<<<<��^���1�uTbJ�k����uz���?Z���������������������<��t��}�)���igt�H���3a�k*������������������������{w2H�j�}M���.2��2к�<<<<<<<<<<<<<<<<<<<<<�9Ӗ�pu����;=dn&��Ak�{��Ż@��r�x�}B�\t�tJ'm:�������s�o�yxxxxxxxxxxxxxxxxxxxx��9S�'���#ө2�VLu��A�_�.К��������������������������^x�DO����s�N�^	�/�Exxxxxxxxxxxxxxxxxxxxx���݀^�=n��C�Nv@S.۝0�%y�X|��<<<<<<<<<<<<<<<<<<<<<��9�I��:ʰ�ɖ~9J��,�%����O�ȼ���������������������� �Y��dec���lv���y�
��zǋ��yxxxxxxxxxxxxxxxxxxxx��݀�fv�z   �?;�z��Sq:�)����^{�A"������������������������� �I�z�vHF���t��,������:q=���<<<<<<<<<<<<<<<<<<<<<�9i`g�z�t@�:�p�z�G��[�k�^�����������������������I&t��D��ge�_O��N�~�F֛/����������������������|��t���Ҟ�޵��OgH����'��,�3<��[�7-�u\�-�#��w�}Mw���������������������|��|����׏I��� �!��n����yxxxxxxxxxxxxxxxxxxxx��9�xu���}���(#��wo|����~���������������������<�s2\ݝ��ki(˿�����Đ��<<<<<<<<<<<<<<<<<<<<<��$tt;|f��;$ש��-˜v��yS����������������������<�sVю��e�z����!�=�=eg�{.�e����������������������<�sr�E3����A����>��<��<<<<<<<<<<<<<<<<<<<<<����}w��<�]�����Y�;���_�7yxxxxxxxxxxxxxxxxxxxx>�sVtt]��w����׮�y�l�x�����������������������y��LN�ݨn�ʟ���!N�l��������������������������<�s�@�t���������{�3�fmLs=[�����g&���������������������|��H��8����;�㮾NKL�����:N����������������������=�[�+�:��m�����ߎ�rw�5ϧ{N�^�z��>-�o���7}�3������������������������<�sVS�����+�:'�O�K띇���������������������ӣ��`Ĭ�����#�w���y��V��3<z   ����'���]��A�4��b���P��˳;�<���:Ӱ�_�S}��S=#������3����������������������<�s�4��n��_V��W�n����>i1�܃�<<<<<<<<<<<<<<<<<<<<<�nx/P�|_=M�ޭ���ϝ?��<�<g�؎(W�������Rs�Dz�xλ3��/��h�i���yw�5�G{��F�]e:�I�^�;:�������K�����������������������鞓B)�!�N�輏��
�^_�r�{NQ��yxxxxxxxxxxxxxxxxxxxx��99�p���s@��L�����w�ws�<<<<<<<<<<<<<<<<<<<<<�𜿙�N�C���k�G�Z��gxN�ә�^y�w�{i����?��\�\���������������������<�s2P�2�#�͠��䉬7CI�Ȋ��w���;�ϧ{N���t���<�{��c�Gb6��� Ͽ#kyxxxxxxxxxxxxxxxxxxxx��99��9� � 1�s��]M�At��4��h�������������������������n{��݉�=k�Zw�|�����h�����������������������Y��'c�I���tгM�^�����=��1К�����������������������'�c�ɂt�_F��6�Y7��Ah��yxxxxxxxxxxxxxxxxxxxx��9�f��c��Ĕ��2�����������������������������y��败�:S�+:�7����萑���g°�T6�3<���d�4�Ԧ�:�>'q]d�e�u7�yxxxxxxxxxxxxxxxxxxxx>�s�-���N��wz��LXu�ְ����w����<<<<<<<<<z   <<<<<<<<<<<<���Ĺ��N�t��;$�)�����Z���������������������<�s�bOb��G�Se��������]�5�3<��=�ݽ�,H��xO_����r��_Ƌ���������������������<����{ܺ�=�>�쀦\�;a:K�t����yxxxxxxxxxxxxxxxxxxxx>�sF���u�a��-�r�:,�Y�K���T�y������������������������"�����(�!���������Y�)���������������������<�����7v:�4���t�S���n��^��DVwӝ��������������������������4��j���|�Y�ѝ�u0�zJ/�#yxxxxxxxxxxxxxxxxxxxx>�s��������u��
�X��~�����������������������������L�,[���ʼ����"�h%��7_�����������������������P���黥=��ki7��ΐv���O@wY�gxN�Q��oZ�긐[G&��F�������������������������h��&��eK���N=�;@$Cګ�~7����������������������<�sf��LwW�niQF����������������������������y��d��;��}��P��=�=�!�yxxxxxxxxxxxxxxxxxxxx��9I��v���1�w2H�S'�[�9���4�����������������������y�笢���V�niw�C�{{��,�\��"���������������������y��䪋fZ{���އ'�i�}*b�~yb�yxxxxxxxxxxxxxxxxxxxx���G�y���_?V���|w�����o���������������������|����.�����y훯]���^�"3�����������������������ϙ���Qݔ�z   ?���C���h�������������������������y��܁ �|�+�ͯ�S���zg�ژ�z���=��a�/�L����������������������D�Y��9q^]c�w��]}���"��k�u�"�G{N��Wu&�������)�����k�O��6��xY}Z��T��o�|g���q���������������������y�符����W�uN<\����;�3<�G����YsW���G���-^k�(ۭ��gx�3VOVw���7��i���~'Xϡ��gw�x���u�ao�"�������zF��W����gv���������������������y��i�2�LS��>����\_��}�b���yxxxxxxxxxxxxxxxxxxxx�9��^�T��z��]�[�	�;$-y�x�:�Q����~W}U[��N��.<<<<<<<<<<<<<<<<<<<<<�wg6�_T_��+�:�����k��������t��`��wtH�_���3:��?�����������������������='�R4Cڝ��yw�V����\���x�u���������������������<�sr��j������6�c�����yxxxxxxxxxxxxxxxxxxxx��93A�v��/��;�:��&�)!<<<<<<<<<<<<<<<<<<<<<����3#���n���O��}ƻ�����������������������y��d��e�G:�iiϛA���Yo����k=�̝�wd�O���I��m�y��@u�Z�,�l���A�G����������������������<�srbgs�AAb��"�)����X�i��1К�����������������������#���N��z   {�:���:K1e�_�&К������������������������/�Oư�ܑ��g�����y�{��c�5�<��N��l�邿��mz�n����2к����������������������<�sz�z�ǰ�Q�)ѯe;�����h�����������������������?�iK�u��WtHo�����!#i��τa��l�gxN��� i�7�M�u4}N����@�n����������������������|��L[:��	�����������a�y'����yxxxxxxxxxxxxxxxxxxxx�9�	�s�	�)���$OwH�S"�Ϳ	����������������������y��LŞ�nk�L��<Z1��7}��@k�gx~7�{6�{�Y�9<����;�z%X�����������������������y��wz`��uG{}:�M�lw�t���:`������������������������|��&I�(�'[��(uXL�����W/<�"��<gEDG��=�P�C���#��%+���/��S���������������������y��w���yo��t�iZO�頧tw�;�z�����;�<'��)�i ՞�����<:�;��`��4�^�G(���������������������|�礁���Y�����u;�n��	�{!�3<'��Y�=�/��y=M�;E��JYo���������������������������wK{�{��nt?�!����<<<<<<<<<<<<<<<<<<<<<�𜎣n�ߴ��q!�8�Lzߍ�5�����������������������ў�M��˖��_?&�z~w�H��W��n�/_/���������������������y����ՙ�������,��#ܽ�z   �w7�������������������������puw�����=�,��3z�{C����������������������<�s�����5��c�d�\�N��,s�i��iL����������������������� �YE;��������.x�X����Y�x�E������������������������Uʹ�w�O�Ӧ�T����<�F���������������������<����)_��w���~��sg����q�����������������������\�Y��]tW����7_�z�=���Ef������������������������39w��)+�/��8	 ���/������������������������ϹA���WΛ_������<��1��l1{�ê_�����������������������󉞳"�s<⼺ƪ�h���:-1E�����8E����n���L\���;7$k�S~;2�ݡ�<<<<<<<<<<<<<<<<<<<<<��9mz����̿�~�����t߻������������������������YM��/��p�x�>�?,�w�gxN�^������׏\��[���Q�[i#<<<<<<<<<<<<<<<<<<<<<���g:����w�o��8O��N��C�/��<<<<<<<<<<<<<<<<<<<<<𜯻�L��~EPO�i��M��p���S��������������������������Y��+
d���~Y}�;\ջ�������|sr���������������������<�s��@��}�4��z��,�?w�HZ�<<<<<<<<<<<<<<<<<<<<<�ub;�\ջ������J͝�]xxxxxxxxxxxxxxxxxxxxx�9��4l⿨���W�u^��ݡ�<<<<<<<<<<<<<<<<<<<<<�9/�w��|'�zU�萾���;�gt.Iϧ{N
�h��;��>��+�z}�˹�9E����z   �������������������y��������2m�?�Z����u���������������������<�s�f�:=�>�_�Gw�u�kM�SBxxxxxxxxxxxxxxxxxxxxx��9�OgFz�I���v����ws�s������������������������@���t��Ҟ7����'��%	#+�zޙ;���<<<<<<<<<<<<<<<<<<<<<��9)ړ��۾��ꎵY��,�+v�<������������������������y������H�<��H�E�St5�ѱ�� �c�5�3<�G���v'F��uj�=�u�bʦ��M�5�3<g_���a'�#��A�6=z=������#��@k�xN�� ��&����f�hO�e�u���������������������y�����v�a��S�_�<v���k�7�1К����������������������4�Ӗ��LY��� O;��CF�nϟ	�^S�<<<<<<<<<<<<<<<<<<<<<��޻�A�oP���h���u�1엁��h����������������������hϙ�t��8����!s3a�Z���N.�Z�����������������������<�s���S:i�I����D6��h����������������������ϙ�=����N�y�b�#�o���w��<<<<<<<<<<<<<<<<<<<<<���n@�lv�³ %rx�=}���w��J�~/���������������������������q���t��r���,��u�⻏����������������������t�M�>�Q�-N���Q���fy/Y�/�^xRE�5�xΊ��&+{;���d��G��KVH��;^d����������������������� ��t7�������Ӵ���AO��vw���{�Y�Mwz   �xNZ�S��@2�=���}gyt�Gw�����i(���P����������������������h�I;s׳����+�c=�v��b_��B�gxN2��l%zt_<+��z��w����0��|Y����������������������C=�����������~:C��_?�eyxxxxxxxxxxxxxxxxxxxx��9Gݲ�ii7��Bnq����k�����������������������=盰��-퟿~L:��� �i�v��_�^����������������������ϙū3�]��EY@/G�{���n����������������������������L7�]K{@Y��g���$�t/���������������������y��$����k0;� �� �N�,oY��&�Әr�������������������������v<G/[ջ��]���1�);��s�.��������������������������.�i�%�z�x�M������y�����������������������y���S����?�X�����Y�������������������������󹞳����
����o�v��{f{ŋ̀7�3<gr:�FuSV��_Vq@f��_�懇���������������������s���}��7��O����y4kc���b��w�U�<3����������������������=gEJ�x�yu�U��w�uZb��ﯭ�q�<<<<<<<<<<<<<<<<<<<<<�9�_ԙ��o�wnH�N��vd��C�yxxxxxxxxxxxxxxxxxxxx>�s��2��e�i�S�~����wǝ�������������������������7�_T_��9�p}jXZ�<<<<<<<<<<<<<<<<<<<<<���^#f�]������x�ͣl��Fxxxxxxxxxxxxxxxxxxxxx����tX=Y�%���r�q���`=�*�_��yxxxxxxxxz   xxxxxxxxxxxx�9_wי������������^_է.Οم�������������������������W�p3M���w��ws}o�I�������������������������y��t�{�R���irw�n�'X������yxxxxxxxxxxxxxxxxxxxx�9��vD��w��]�Um��; һ���������������������<�sޝi��Q}ES�L뼖ϻC�yxxxxxxxxxxxxxxxxxxxx>�s^6��*��N�����!}]�w���\���O��J�iw�G�}��WX��ڗs�s��=�������������������������9��5���:d������������������������������y����uz�}b�Џ�X�<�ךx�����������������������<�sҟΌ�ʓ���Ks?�����皇��������������������������p��=o=O'Od�JFV���3w�ߑ-xxxxxxxxxxxxxxxxxxxxx>�sR�'���}�I��k=��YNW�y�Y��������������������������͑y����\��j��c��A��@k�gxN�Xw�;�N��Y�Ժ{��,ŔM��@k�gx�:�0?�NrG֧��mz�z~���IG����<<<<<<<<<<<<<<<<<<<<<��;A�M��2"���ͺў��@�.������������������������5���^G%�D��y�L_�מo�c�5�3<�h@�-�י�^�!�A�v�G���ݞ?����yxxxxxxxxxxxxxxxxxxxx��9�w'��ޠ6����9��"c�/�������������������������ў3m�W'p��/��C�fª����\���/���������������������y���'$�E'L�tҦ�<�! 9N1�l<z   7�&К����������������������3{��=2�*�h�TG�������yxxxxxxxxxxxxxxxxxxxx���݀����gAJ���{�:0���`�2^�������������������������5�����1��d4�2��	�Y����w�����������������������3�$}��[�l闣�9`1��^��_\���k<<<<<<<<<<<<<<<<<<<<<�MV�0v@I�fw�<�����w��:N�������������������������nf���ө�i=�������p���$����<<<<<<<<<<<<<<<<<<<<<𜴮�h��dT{�O����蘏���Pza�����������������������ў�v�gMT�#W��z���ž&��<<<<<<<<<<<<<<<<<<<<<��dBg�J��xV���4��G+ad���>χzN'O�-���]K���t���/�~�����������������������<�s:��e��nPǅ��82�}7��t7�G{�7a/[�?��t���"�^����|������������������������3�Wg���wK��2��^�p��w����7�3<'��ݙn���������I	�^�����������������������IBG���`v�A��Ar�:Y޲�i�M��1�>�<g�x�^��wK���b�c�Svf���]	�3<'W]4��K��><�N��S���������������������������?�w�|�c������ϝ廳����}����������������������s=gEGw�\}W�k�|�������o�gx��t܍ꦬ�鿬�$��F��/��z   3<�I��^9o~���_��;�h��4׳�,����~yf"�'zΊ��������=������_[��yxxxxxxxxxxxxxxxxxxxx>�s��"�3q��V�ܐ��N���,w�^���������������������|���e�����2����~��;�}�;�3<g5�o�­s��������yxxxxxxxxxxxxxxxxxxxx��9=z�F̚���_?r}Wo�Z�G�n�����������������������<��	�z��K�տ�N�<-�;�zUL�<����������������������<�s��3{�A=է�7�3½��O]�?��3<gMS�(��f��e�9�pU�������=����������������������� ������������JO�H���#i����������������������<�s�1��rU������*5w:@�w���������������������y��;Ӱ������^��y-�w�^���������������������|��l��U���U��C���N�<�ѹ$�1<<<<<<<<<<<<<<<<<<<<<��9)������������/���{�������������������������sWk<?�tȴ��k}7��������������������������	����0�~�ݱ�y4�5�N	���������������������y��?��'}w���~�m��3��u�5�3<'�/�?��NK{�z�N��z3�$��X�yg�̿#[���������������������|��hOJwo�Γ��;�zd!f������;�������������������������3;�#�#=�N��DD�ZO�����<<<<<<<<<<<<<<<<<<<<<����w؝ݳ֩u���Y�)���7��<<<<<<<<<<<<<<<<<<<<z   <��u|a~2��䎬O=�����N�;ߓ���yxxxxxxxxxxxxxxxxxxxx�9�w�<f�,H�eDHoӛu�=����]������������������������k��=���JL�~-�ؙ�N�=���@k�gx�рN[��3e��Cz�<��I�=&{Me���������������������<�sz�NI#�Am����s�Eư_Zw�����������������������=g���N�t_x���̈́U7h{�;�xh�_���������������������� ϹOH��N�N�M'y�C@r�b�xn�M�5�3<g*�$v[{d:U�ъ����!����Z���������������������<��ݳ��ς�����u>`��)�+��e��3<��k �ǭ;�c���h�e`���$O���>�����������������������=g4I�XG�8��/G�s�b��d��z�I��xxxxxxxxxxxxxxxxxxxxx�9+":���a쀒���y>/Y!�_�x�u�"�<�����{�g�SO�z*N=������k��/Hdu7�yxxxxxxxxxxxxxxxxxxxx�9i]O�Nɨ�ܟ�����1�Y_#�����>B����������������������='��]Ϛ�^G�P�����w�}M��yxxxxxxxxxxxxxxxxxxxx��9Ʉβ���}����i�)ҏV��z�e}���N��[ڳ߻�v���iw_|�t����������������������y��tu����ݠ���qd��n���n����o�>^����1���D2����w#|�z!�3<g��tw���ed�������o�gxN���3��wz   -�e�7�ѳߓн��������������������������n�����x'��:u��e��N�<Oc�}�x�*���lU�vw�;ĺǰ���r�Ż,�gxN��h����;�}x�6ݧ"���!6�����������������������4��N��Ǿ����cU�;�wg]����&��zΊ��+����׾���;��/2�<<<<<<<<<<<<<<<<<<<<<�����MY��Y=�I ����_��gx�����r��Z?տ~�w�Ѭ�i�g�Y؃�V���D�O��)����5V}G{���i�)r���^�)���������������������|��t|EPg����޹!Y;��ۑY������������������������t�i��P��էe�M�����w���w�gx�j���Q}�[������ai����������������������<�sz�z��5w���~�����6���J���������������������y��?�a�du���3ȝ�yZ�w����~yv���������������������y��|�]g��+�z�O;�o�g�{}U��8f�gxΚ�^Q ��4���s�����5��'-�{��������������������������J�﫧��ջ��`����GҒ���������������������y��c�����w�W�Uj�t�H����������������������� �yw�a�E�M�2��Z>������������������������h�y���L�;	֫zG���u��y>�sI�cxxxxxxxxxxxxxxxxxxxxx>�sR(E3��I��qW_a��k_�u�)��\7�3<'���x~���i��z   1��.�n�������������������������7��a�a��B?�c��h^k������������������������I:3�+O��v/������g���k�gxN�_f�Ý����<�<��f(IY����ܙG�����������������������t�Iў�����'}Tw���B�f9]���wd-�3<'g v6G�$Fz.r����>������yxxxxxxxxxxxxxxxxxxxx��9=b�m�4�;1�g�S��S6��o�yxxxxxxxxxxxxxxxxxxxx��9����d;�Y�z�������w�'�?Z���������������������<�s��y�6Y�.�ˈ�ަ7�F{:�/��8�3<�׬�{{���Z�3}�^{�Ꮑ�<<<<<<<<<<<<<<<<<<<<<������t_g�zE��y��2�v{�L������������������������y���ޝ�Fx��t_G��$���a���F;�G{δ�3\���>��N��	�n���wr�.к������������������������s��8�0��I�N�t���8� �����@k�gx�T�I���t�̣SqC��������������������������y��w�g���)�����|�ܿS�W���x�gx~7�� v�[w��Ч�Д��v'LgI���}<ϧ{�h����2lq��_�R��4�{�:~q�*2����������������������<�sVDt4Y���%=$��=�|^�B����"�8E�x~7�������N����T�zJw��í���_���n����������������������<�sҺ����Q�?��;ˣc>���Fz   \OC�}�"�G{Nؙ��5P��8\��Q����� ����������������������<�s�	�e+ѣ��Y����4�S��������<<<<<<<<<<<<<<<<<<<<<�9�<}��g�w-�F������	�.������������������������8��MK�Ar��Ȥ��h_��<<<<<<<<<<<<<<<<<<<<<�9߄}�li���cҩ�w�dH{���F���B�gx�,^���j�-�/��z9���}�w��<<<<<<<<<<<<<<<<<<<<<��Wwg���Z���o>�g�'1$�{!�3<'	�_��9�N�u�dy�2��6y�Ɣ�<<<<<<<<<<<<<<<<<<<<<�U��9z٪�-��w�u�aOٙ型wY$<<<<<<<<<<<<<<<<<<<<<��\u�Lk/qw����;m�OE��/�Cl4�3<�h@ߝ�5�}W���Ǫ>w��κ���M�����EWp�]=�}�w�3�+^d�yxxxxxxxxxxxxxxxxxxxx��9��q7������z�� 2��B�0?<<<<<<<<<<<<<<<<<<<<<��;$��{���~��^�̣Y�\����;��噉<<<<<<<<<<<<<<<<<<<<<��9+R:�#Ϋk��������S�~m��S����������������������h��������[�sC�v:�#��z�����������������������Ӧ��/�O������M��L��;�<<<<<<<<<<<<<<<<<<<<<��������
�Ή��S���z���������������������y�����:1k��?���]��kme��6�����������������������&�����.qW�f�;�����9T1������������������������� �����4��W�T�v��T����>z   uq��.<<<<<<<<<<<<<<<<<<<<<��5M��@��i����U���kx�OZ�7� 7�<���*�WO���w+=�"�s珤%���������������������� �Y� �#�U���絛j���� �ޅ������������������������L�&���+�zeZ�|�z����������������������ў�~W��w�W�����:��|F������������������������|��P�fH��>:�㮾ª�׾��S�n�gxN�1\�����! �&�c��]��\7�3<�o&�������~t�Z�Ѽ��;%�������������������������tf�W����^��i����x7�=�<<<<<<<<<<<<<<<<<<<<<��T���H�;-�y3�y:y"��P�0�b�睹3��l����������������������鞓�=)ݽ�;O���X둅��r�b7����Z�gxN�@�l�4�#H��\�:EW}k=�?Z���������������������<�szĺ��i`wbt�Z���#_g)�l���Z���������������������<�s����v�;�>�lӣ��;=�|O:�����������������������y����	�m� ]�!�Mo֍�t�_Zwq�gxN�Yo��:*1%���cg�:��|��yxxxxxxxxxxxxxxxxxxxx���G:m�Δ����?:d$����0�5�������������������������;$���龎��I\�~hݍv����;ʍI� Zg�|�s���-k毉E�����HD������������|��L[:��	�����������a�y'��{�<<<<<<<<<<<<<<<<<<<<<���Ĺ��N�t��;$�)z   ����Z���������������������<�s�bOb��G�Se���{A�;h����������������������ϟt�fw/<R"�'�����ܿS�W���x�gx�4�� v�[w��Ч�Д��v'LgI���m�����������������������=g4I�XG�8��/G�s�b��d��z�I��xxxxxxxxxxxxxxxxxxxxx�9+":���a쀒���=�l/Y!�_�x�u�"�<����{�g�SO�z*N=���������_���n����������������������<�sҺ����Q�?��;ˣc>���F\OC�}�"�G{Nؙ��5P��8\��Q����� ����������������������<�s�	�e+ѣ��Y����4�S��������<<<<<<<<<<<<<<<<<<<<<�9�<}���{�Zڍ�3��}���]������������������������q�-�NK�Ar��Ȥ��h_��<<<<<<<<<<<<<<<<<<<<<�9_�}�li���cҩ�w�dH{���F���B�gx�,^���j�-�ߔ��r��?|����~���������������������<�s2\ݝ��ki(˿�F�~ObH@�B�gxN:���s������eN;m�<�)�yxxxxxxxxxxxxxxxxxxxx�9�h�s��U�[����Þ�3�=�Hxxxxxxxxxxxxxxxxxxxxx��9�ꢙ�^����w�t��ؿ_���h�gx�р�;�k����׏U}�,ߝu}�/�<<<<<<<<<<<<<<<<<<<<<��9+:�����z^�b��w�3�+^d�yxxxxxxxxxxxxxxxxxxxx��9��q7����Y=�I ���B�0?<<<<<<<<<<<<<<<<<<z   <<<��;$��{��{�T��{�3�fmLs=���=��a�/�L����������������������D�Y��9q^]c�w��]}���"�����8E����n���L\������)�����k�O��6��xY}Z�_T��o��3������������������������<�sVS�����+�:'�����z���������������������y�����:1k��?���]��km�s+m������������������������O@�Փ�]��� w�i��	�s�b���:�<���u�a~EPO�i��zF�׮����3_���������������������y��i�2�LS��>����\_��}�b�܃�<<<<<<<<<<<<<<<<<<<<<�nx/P�|]=M�ޭ���ϝ?��<�<g�؎(W�������Rs�D�+<<<<<<<<<<<<<<<<<<<<<�wg6�?T_��+�:�e{w�5�G{��F�]e:�I�^�;:����γ��%�����������������������|��P�fH��>:�㮾ª�n_�u�)��\7�3<'���x~�tȴ��k}7��������������������������uz�}b�Џ�X�<�ךx�����������������������<�sҟΌ�ʓ���Ks?����ws�s������������������������@���t��Ҟ7����'��%	#+�zޙ;���'xxxxxxxxxxxxxxxxxxxxx>�sR�'���}�I��k=�󱜮���;�������������������������3;�#�#=�N��DD�ZO�����<<<<<<<<<<<<<<<<<<<<<����w؝ݳ֩u���Y�)�����<<<<<<<<<<<<<<<<<z   <<<<��u|a~2��䎬O=�������w����_�yxxxxxxxxxxxxxxxxxxxx�9�w�<�3Y�.�ˈ��L��頿���<<<<<<<<<<<<<<<<<<<<<��^���1�uTbJ�k����uz���_�yxxxxxxxxxxxxxxxxxxxx���G:m�Δ����igt�H���3a�k*��������������������������d�4�Ԧ�:�>'q]d�e�u7�yxxxxxxxxxxxxxxxxxxxx>�s�-���N��wz��LXu�ְ����w�ֽs�x�}B�\t�tJ'm:�����ȇ��w�yxxxxxxxxxxxxxxxxxxxx��9S�'���#ө2�VLuĽ������������������������y��O�g���)�����l`��)�+��e��3<�k �ǭ;�c���h�e`���$O���6�����������������������3�$}��[�l闣�9`1��^��_\���k<<<<<<<<<<<<<<<<<<<<<�MV�0v@I���y�����w��:N�����������������������?�nf���ө�i=�������p����/Hdu7�yxxxxxxxxxxxxxxxxxxxx�9i]O�Nɨ�ܟ�����1�Y_#�����>B����������������������='��]Ϛ�^G�P�����w�}M��yxxxxxxxxxxxxxxxxxxxx��9Ʉβ���}����i�)ҏV��z�e}���N��[��w-�F������	�.������������������������8�}��ݠ���qd��n���n����/�>^����1���D2����w#|�z!�3<g��tw���o��z9������f�yxxxxxxxxxxxxxxxxxxxx��9���z   tsߵ���_l�g�'1$�{!�3<'	�_��9�N�u�dy�2��6y�Ɣ�<<<<<<<<<<<<<<<<<<<<<�U��9z٪�-��w�u�aOٙ型wY$<<<<<<<<<<<<<<<<<<<<<��\u�Lk/qw����;m�OE��/�Cl4�3<�h@ߝ�5�}W���Ǫ>w��κ���M�����EWp�]=�}���;��/2�<<<<<<<<<<<<<<<<<<<<<�����MY��߬�$�̇��_��gx�����r���~����ޙG�6���O�����g&���������������������|��H��8����;�㮾NKL�����u�"�G{N��Wu&��m�����ߎ�rw�5ϧ{N�^�z��>-�/���7}���{w�yxxxxxxxxxxxxxxxxxxxx��9�)~s�C�n��V{ci����������������������<�sz�z��5w���~�����6��6������������������������'�����.qW�b�;�����9T1��|��������������������������:Ӱ?�"����ÿS=#�kW}��������������������������<�s�4��n��_V��W�n����>i1{�An�xN7�(U���&wW�Vz�E���IK�������������������������AlG��z���U_�V���"��xλ3����h�i�ײ�;�����������������������=�e#��2��$X�����uz��F��fxxxxxxxxxxxxxxxxxxxxx>�sR(E3��I��qW_a�k�/���{�������������������������sWk<?�:dz   ������������������������������y��|g�:=�>�_�Gw�u�kM�SBxxxxxxxxxxxxxxxxxxxxx��9�OgFz�I���v���ƻ�����������������������y��d��e�G:�iiϛA���Yo����k=�̝�w�<<<<<<<<<<<<<<<<<<<<<��9)ړ��۾��ꎵY��XNW�y�Y��������������������������͑y����\��j��c��A��@k�gxN�Xw�;�N��Y�Ժ{��,ŔM��@k�gx�:�0?�NrG֧�������N�;�IG����<<<<<<<<<<<<<<<<<<<<<��;A�,H�eDH�?֍�t�_Zwq�gxN�Yo��:*1%���cg�:���ᯁ�<<<<<<<<<<<<<<<<<<<<<������t_g�zE���?:d$����0�5�������������������������ow2H�j�}M���.2��2к�<<<<<<<<<<<<<<<<<<<<<�9Ӗ�pu����;=dn&��Ak�{��Ż@��9�<�>!q.:a:��6����q�A��s�;��<<<<<<<<<<<<<<<<<<<<<��ؓ�m��T�G+�:��C����Z���������������������<��ݳ��ς�����u60���`�2^�����������������������?�5�����1��d4�2��	�Y����w�����������������������t�M�>�Q�-N���Q���fy/Y�/�^xRE�5�xΊ��&+{;����cw�<�KVH��;^d����������������������� ϟt7�������Ӵ���AO��vw�����$����<<<<<<<<<<<<<<<<<<<<<𜴮�h��dT{�O����蘏�z   ����Pza�����������������������ў�v�gMT�#W��z���ž&��<<<<<<<<<<<<<<<<<<<<<��dBg�J��xV���4��G+ad���>χzN'O�-��޻�v���iw_|�t����������������������y��tu˾��nPǅ��82�}7��t7�G{�a/[�?��t���"�^����|������������������������3�Wg���wK�7ed����}�w��<<<<<<<<<<<<<<<<<<<<<��Wwg���Z���/�ѳߓн��������������������������n�����x'��:u��e��N�<Oc�}�x�*���lU�vw�;ĺǰ���r�Ż,�gxN��h����;�}x�6ݧ"���!6�����������������������4��N��Ǿ����cU�;�wg]����&��zΊ��+����׾��������o�gx��t܍ꦬ��oVq@�C��/��3<�I��^9o�^?��^�̣Y�\�'fa~wX��3yxxxxxxxxxxxxxxxxxxxx>�sV�t�G�W�X��qW_�%������:N����������������������=�[�+�:���z�d�t�oGf�;������������������������=�M/C=^V�������>�L��;�<<<<<<<<<<<<<<<<<<<<<��������
�Ή�k�����yxxxxxxxxxxxxxxxxxxxx��9=z�F̚���_?r}Wo�Z�G��J���������������������y����a�du���1ȝ�yZ�w����~y����������������������� ��}w�i؟_�S}��ߩ��z   ��>uq��Wxxxxxxxxxxxxxxxxxxxxx��9k�zE�7��/��q��z7���v���=� 7�<���*_WO���w+=�"�s珤%���������������������� �Y� �#�U���絛j���� ��
�<�ݙ�M��W4�ʴ�k��z����������������������ў�~W��w�W�����:��l�sIz3<<<<<<<<<<<<<<<<<<<<<��9)����������ۗs�s��=�������������������������9��5��{2m��Z����u���������������������<�s�3A�v��/��;�:��&�)!<<<<<<<<<<<<<<<<<<<<<����3#���n���O��}o��\�\���������������������<�s2P�2�#�͠��䉬7CI�Ȋ��w���;�	�O���I��m�y��@u�Z�,�|,�+v�<������������������������y������H�<��H�E�St5�ѱ�� �k�5�3<�G���v'F��uj�=�u�bʦ��E�5�3<g_���a'�#��A�gz�z~����#��@k�xN�� ��L��2"�?��F{:�/��8�3<�׬�{{���Z�3}�^{���@k�gx�рN[��3e��C�y��2�v{�L������������������������y����;$���龎��I\�~hݍv����iKg�:��}|�27Vݠ5�=���]�u���������������������s��8�0��I�N�t���8� ����@k�gx�T�I�z   ��t�̣Sq�!�{���yxxxxxxxxxxxxxxxxxxxx���Ӏ����gAJ���{�:��w��J�~/����������������������ϟ���q���t��r���,��u������������������������|��&I�(�'[��(uXL�����W/<�"��<gEDG��=�P�C�G��%+���/��S���������������������y��O���yo��t�iZO�頧tw�;�z}{�Y�Mw�xNZ�S��@2�=���}gyt�Gw�����i(���P����������������������h�I;s׳����+�c=�v��b_��B�gxN2��l%zt_<+��z��w����0��|Y����������������������C=�����|�]K���t���/�~�����������������������<�s:��e�ii7��Bnq����k�����������������������=狰��-퟿~L:��� �i�v��_�^����������������������ϙū3�]���2��^�p������o�gxN���3��w-�e�����I	�^�����������������������IBG���`v�A��Ar�:Y޲�i�M��1�>�<g�x�^��wK���b�c�Svf���]	�3<'W]4��K��><�N��S���������������������������?�w�|�c������ϝ廳����}����������������������s=gEGw�\}W�k_�v��{f{ŋ̀7�3<gr:�FuSV��7��8	 ��_�懇���������������������s���}��7����w�Ѭ�i�����;��z   噉<<<<<<<<<<<<<<<<<<<<<��9+R:�#Ϋk��������S�~}z�����������������������ў�-�A���[�sC�v:�#��z�����������������������Ӧ��/�O������M�}���w�gx�j����P}�[��õ��XZ�<<<<<<<<<<<<<<<<<<<<<���^#f�]������x�ͣ|n�����������������������<���	�z��K�տ�N�<-�;�zUL�<_���������������������y������4�ϯ�>���T���U��8�+<<<<<<<<<<<<<<<<<<<<<��5M��@��i����U���kx�OZ̞{��������������������������J������ջ��`����GҒ���������������������y��c�����w�W�Uj�t�H�������������������������L�&���+�zeZ�l������������������������h�y���L�;	֫zG���u��y�ѹ$��O��J�iw�G�}��WX���˹�9E�����������������������y������Ͻ��6�_c�����yxxxxxxxxxxxxxxxxxxxx��9ߙ�N�C���k�G�Z��gxN�ә�^y�w�{i������n�{�yxxxxxxxxxxxxxxxxxxxx��9�~���wZ��f��t�D֛�$ad�Z�;sg��ϧ{N���t���<�{��c�Gb>���A�G����������������������<�srbgs�AAb��"�)����X�i��5К�����������������������#���N��{�:���:K1e�_�"К������������������������/�Oư�ܑ���3=z=����~��k�5z   �<��N��|&�ҟ�u�=�����S�  :_IDAT�]������������������������k��=���JL�~-�ؙ�N�={�k�5�3<�h@�-�י�^�!��<��I�=&{Me���������������������<�s�۝�Fx��t_G��$���a���F;�G{δ�3\���>��N��	�n���wr�.кw���������������������� ϹOH��N�N�M'y�C@r�b����N�5�3<g*�$v[{d:U�ъ�������w��<<<<<<<<<<<<<<<<<<<<<���i@�lv�³ %rx�=}���;�z%X�����������������������y��Oz`��uG{}:�M�lw�t���:`���yxxxxxxxxxxxxxxxxxxxx>�sF���u�a��-�r�:,�Y�K���T�y������������������������"�����(�!���#�������Y�)���������������������<�����7v:�4���t�S���n�������;�<'��)�i ՞�����<:�;��`��4�^�G(���������������������|�礁���Y�����u;�n��	�{!�3<'��Y�=�/��y=M�;E��JYo���������������������������wK{������~:C��_?�eyxxxxxxxxxxxxxxxxxxxx��9Gݲﴴ�q!�8�Lzߍ�5�����������������������ў�E��˖��_?&�z~w�H��W��n�/_/���������������������y����ՙ�����MY@/G���w����7�3<'��ݙn�����m���$�t/�������z   ��������������y��$����k0;� �� �N�,oY��&�Әr�������������������������v<G/[ջ��]���1�);��s�.��������������������������.�i�%�z�x�M������y�����������������������y���S����?�X�����Y�������������������������󹞳����
����/v�z�=���Ef������������������������39w��)+���C�����/������������������������ϹA���WΛ��O�߿�;�h��4��Y؃�V���D�O��)����5V}G{���i�)r��>��S����������������������h����������޹!Y;��ۑY������������������������t�i��P��էe�E�����>�}�;�3<g5�o���­s���jo,�w�gxN�^������׏\��[���Q>��Fxxxxxxxxxxxxxxxxxxxxx����tX=Y�%��_r�q���`=�*�_�����������������������<�s~�]g��W�T�v�w�g�{�O]�?��gxΚ�^Q ��4���s�����5��'-f�=����������������������� ������������JO�H���#i����������������������<�s�1��rU������*5w:@������������������������ �yw�a�C�M�2��Z�w�^���������������������|��l��U���U��C���N�<��\��ϧ{N
�h��;��>��+�z���\���x�u���������������������<�sr��j����@��L�����w�ws�<<<<<<<<<<<<<<<z   <<<<<<���LP��݇!��莵Σy��wJ�3<'���H�<�۽4��n{��x7�=�<<<<<<<<<<<<<<<<<<<<<��T���H�;-�y3�y:y"��P�0�b�睹3��|�����������������������='E{R�{�w��=Pݱ�#1��� Ͽ#kyxxxxxxxxxxxxxxxxxxxx��99��9� � 1�s��]M�At��4��h�������������������������n{��݉�=k�Zw�|�����h�����������������������Y��'c�I���t������yg?��5К�����������������������'�c>�邿����Ǻў��@�.������������������������5���^G%�D��y�L_�מ=�5К����������������������4�Ӗ��LY���@�v�G���ݞ?����yxxxxxxxxxxxxxxxxxxxx��9��NI#�Am����s�Eư_Zw�����������������������=g���N�t_x���̈́U7h{�;�xh�;���������������������y���'$�E'L�tҦ�<�! 9N1�|xn~'К����������������������3{��=2�*�h�TG�{����@k�gx�4�{6�{�Y�9<�����r��_Ƌ���������������������<����{ܺ�=�>�쀦\�;a:K�t��n�<<<<<<<<<<<<<<<<<<<<<��9�I��:ʰ�ɖ~9J��,�%����O�ȼ���������������������� �Y��dec���|��g{�
��zǋ��yxxxxxxxxxxxxxxxxxxxx��Ӏ�fvޛ?;�z��Sq:�)����^�^��DVwӝ��������������������������4��j���|�Y�ѝ�u0�zJ/�#yxxxxxxxxxxxxxxz   xxxxxx>�s��������u��
�X��~�����������������������������L�,[���ʼ����"�h%��7_�����������������������P���黥=�{��nt?�!����<<<<<<<<<<<<<<<<<<<<<�𜎣n�wZ�긐[G&��F�������������������������h��"��eK���N=�;@$Cګ�~7����������������������<�sf��LwW�ni���,��#�����n����������������������������L7�]K{@Y��6z�{C����������������������<�s�����5��c�d�\�N��,s�i��iL����������������������� �YE;��������.x�X����Y�x�E������������������������Uʹ�w�O�Ӧ�T����<�F���������������������<����)_��w���~��sg����q�����������������������\�Y��]tW�����]���^�"3�����������������������ϙ���Qݔ�?���!N�|h�������������������������y��܁ �|�+��������y4kc����,����~yf"�'zΊ��������=������_�^�)���������������������|��t|EPg���V�ܐ��N���,w�^���������������������|���e�����2����~�g��wǝ�������������������������7�?T_��9�pm�7��;�3<�G����YsW���G���-^k�(�[i#<<<<<<<<<<<<<<<<<<<<<���:����w�/��8O��N��C�/��yxxxxxxxxxxxxxxxxxxxx�9��3��+�z�O;�;�3½vէ.Ο�
z   �3<gMS�(��f��e�9�pU�����������������������������y��t�{�R���irw�n�'X������yxxxxxxxxxxxxxxxxxxxx�9��vD��w��]�Um��; �_���������������������y��;Ӱ������^��y-ۻC�yxxxxxxxxxxxxxxxxxxxx>�s^6��*��N�����!}]�w�mt.Io�����������������������='�R4Cڝ��yw�V�v�r�{NQ��yxxxxxxxxxxxxxxxxxxxx��99�p���so�C@�M��X����n�gx�w&�������~t�Z�Ѽ��;%�������������������������tf�W����^��i���m���k�gxN�_f�Ý����<�<��f(IY����ܙG>����������������������鞓�=)ݽ�;O���X둅���t�n��ߑ�<<<<<<<<<<<<<<<<<<<<<�𜜁��i�G���u��&� :�z�����������������������y���u������螵N��G��RL��׿����������������������y����1�$wd}:��L�^������t��h���������������������� ���1�ɂt�_F��g�c�hO�e�u���������������������y�����v�a��S�_�<v���k��h�����������������������?�iK�u��WtH O;��CF�nϟ	�^S�<<<<<<<<<<<<<<<<<<<<<���v'��ޠ6����9��"c�/�������������������������ў3m�W'p��/��C�fª����\������������������������<�s���S:i�I����D><7�h����������������������ϙ�=����N�y�b�#�=}��]�5z   �3<�=�ݽ�,H��xO_gs�N�^	�/�Exxxxxxxxxxxxxxxxxxxxx���Ӏ^�=n��C�Nv@S.۝0�%y�X|�y�O���$�ce��dK����i���u���'Ud^���������������������y�笈�h����JzH>v�ȳ�d�t��E�q�<<<<<<<<<<<<<<<<<<<<<��i@w3;�͟�N=M�8���nw�[�o�A"������������������������� �I�z�vHF���t��,������:q=���<<<<<<<<<<<<<<<<<<<<<�9i`g�z�t@�:�p�z�G��[�k�^�����������������������I&t��D��ge�_O��N�~�F֛/����������������������|��t���Ҟ�ki7��ΐv���O@wY�gxN�Q��;-�u\�-�#��w�}Mw���������������������|��|����׏I��� �!��n����yxxxxxxxxxxxxxxxxxxxx��9�xu���}��SF������w7�������������������������puw�����=�,�b=�=�!�yxxxxxxxxxxxxxxxxxxxx��9I��v���1�w2H�S'�[�9���4�����������������������y�笢���V�niw�C�{{��,�\��"���������������������y��䪋fZ{���އ'�i�}*b�~yb�yxxxxxxxxxxxxxxxxxxxx���G�y���_?V���|w�����o���������������������|����.�����y�ݮ�y�l�x�����������������������y��LN�ݨn�ʟ�f�'d>��������������������������<�s�@�t������S�����<��1��|b��w�U�<3����������������������z   =gEJ�x�yu�U��w�uZb���O��yxxxxxxxxxxxxxxxxxxxx>�s��"�3q�o�wnH�N��vd��C�yxxxxxxxxxxxxxxxxxxxx>�s��2��e�i�Q�~���t߻������������������������YM����p�x���K띇���������������������ӣ��`Ĭ�����#�w���y�ϭ��gx�?VOVw�����i���~'Xϡ����<<<<<<<<<<<<<<<<<<<<<��wי���A=է����^��S��|��������������������������W�p3M���w��ws}o�I��sr���������������������<�s��@��u�4��z��,�?w�HZ�<<<<<<<<<<<<<<<<<<<<<�ub;�\ջ������J͝����������������������<�sޝi���P}ES�L뼖�ݡ�<<<<<<<<<<<<<<<<<<<<<�9/�w��|'�zU�萾���;�6:��7����������������������鞓B)�!�N�輏��
�^�}9�=�(�s�<<<<<<<<<<<<<<<<<<<<<��c�Z���7�! �&�k��]��\7�3<�;��a�a��B?�c��h^k������������������������I:3�+O��v/������6��u�5�3<'�/�?��NK{�z�N��z3�$��X�yg�̿#�����������������������t�Iў�����'}Tw���B��r�b7����Z�gxN�@�l�4�#H��\�:EW}k=�Z���������������������<�szĺ��i`wbt�Z���#_g)�l��_Z���������������������<�s����v�;�>�|�G��wz��O:�����������������������y����	�z   ��dA��/#B�3��n����2к����������������������<�sz�z�ǰ�Q�)ѯe;���g����������������������y��败�:S�+:�?�����!#i��τa��l�gxN��A�oP���h���u�1엁��h����������������������hϙ�t��8����!s3a�Z���N.�Z��yxxxxxxxxxxxxxxxxxxxx�9�	�s�	�)���$OwH�S"���	����������������������y��LŞ�nk�L��<Z1����w�.К����������������������?���^x�DO�������\���"<<<<<<<<<<<<<<<<<<<<<���i@����h��O';�)���N�Β<],��<ϧ{�h����2lq��_�R��4�{�:~q�*2����������������������<�sVDt4Y���%=$�{��^�B����"�8E�x�4�������N����T�zJw��í׷׿ ���t���������������������y��u=E;$��s:�w�G�|tg}������E����4�3w=k:�zq�B=֣n��-�5~/���������������������y��$:�V�G�ų2ﯧix�H?Z	#�͗�yxxxxxxxxxxxxxxxxxxxx>�s:y�ni��޵��OgH����'��,�3<��[���v�:.�ǑI�Ѿ��yxxxxxxxxxxxxxxxxxxxx>�s��x�����ǤS��ɐ�j�ߍ���<<<<<<<<<<<<<<<<<<<<<��Y�:��վ[ڿ)#��w������������������������y��d��;��}��P������Đ��<<<<<<<<<<<<<<<<<<<<<��$tt;|f��;$ש��-˜z   v��yS����������������������<�sVю��e�z����!�=�=eg�{.�e����������������������<�sr�E3����A����>��<��<<<<<<<<<<<<<<<<<<<<<����}w��<�]�����Y�;���_�7yxxxxxxxxxxxxxxxxxxxx>�sVtt]��w����nW�g�W��x���������������������<�s&��nT7e�O�z�� 2Z��~a~xxxxxxxxxxxxxxxxxxxxx��9w H:���y�������zg�ژ�z>1{�ê_�����������������������󉞳"�s<⼺ƪ�h���:-1E��ק�q�<<<<<<<<<<<<<<<<<<<<<�9�_ԙ����;7$k�S~;2�ݡ�<<<<<<<<<<<<<<<<<<<<<��9mz����̿�~����g���q���������������������y�符����W�uN<\[퍥���������������������������u0b�������z���<��V��3<����'���]��A�4��b���P����u�x���L���������N��p�]����g������������������������Y��+
d���~Y}�;\ջ���������yxxxxxxxxxxxxxxxxxxxx�9��^�T��z��]�[�	�;$-y�x�:�Q����~W}U[��N��Wxxxxxxxxxxxxxxxxxxxxx�9��4l�����W�u^����k��������t��`��wtH�_��g�Kқ����������������������t�I�͐v'}t��]}�U�ݾ��S�n�gxN�1\������i��5��.�n�������������������������	����0�~�ݱ�y4�5�N	�������z   ��������������y��?��'}w���~�m�{��皇��������������������������p��=o=O'Od�JFV���3w�ߑO���������������������|��hOJwo�Γ��;�zd!�c9]���wd-�3<'g v6G�$Fz.r����>�����_�yxxxxxxxxxxxxxxxxxxxx��9=b�m�4�;1�g�S��S6��/�yxxxxxxxxxxxxxxxxxxxx��9����d;�Y�z>ӣ��;=��'�Z���������������������<�s��y�g� ]�!���X7��Ah��yxxxxxxxxxxxxxxxxxxxx��9�f��c��Ĕ��2�����ڳ��Z���������������������<��t��}�)������萑���g°�T6�3<���� i�7�M�u4}N����@�n����������������������|��L[:��	�����������a�y'��{�<<<<<<<<<<<<<<<<<<<<<���Ĺ��N�t��;$�)����Z���������������������<�s�bOb��G�Se���{A�;h����������������������ϟt�fw/<R"�'�����ܿS�W���x�gx�4�� v�[w��Ч�Д��v'LgI���m�����������������������=g4I�XG�8��/G�s�b��d��z�I��xxxxxxxxxxxxxxxxxxxxx�9+":���a쀒���=�l/Y!�_�x�u�"�<����{�g�SO�z*N=���������_���n����������������������<�sҺ����Q�?��;ˣc>���F\OC�}�"�G{Nؙ��5P��8\��Q����� ����z   ������������������<�s�	�e+ѣ��Y����4�S��������<<<<<<<<<<<<<<<<<<<<<�9�<}���{�Zڍ�3��}���]������������������������q�-�NK�Ar��Ȥ��h_��<<<<<<<<<<<<<<<<<<<<<�9_�}�li���cҩ�w�dH{���F���B�gx�,^���j�-�ߔ��r��?|����~���������������������<�s2\ݝ��ki(˿�F�~ObH@�B�gxN:���s������eN;m�<�)�yxxxxxxxxxxxxxxxxxxxx�9�h�s��U�[����Þ�3�=�Hxxxxxxxxxxxxxxxxxxxxx��9�ꢙ�^����w�t��ؿ_���h�gx�р�;�k����׏U}�,ߝu}�/�<<<<<<<<<<<<<<<<<<<<<��9+:�����z^�b��w�3�+^d�yxxxxxxxxxxxxxxxxxxxx��9��q7����Y=�I ���B�0?<<<<<<<<<<<<<<<<<<<<<��;$��{��{�T��{�3�fmLs=���=��a�/�L����������������������D�Y��9q^]c�w��]}���"�����8E����n���L\������)�����k�O��6��xY}Z�_T��o��3������������������������<�sVS�����+�:'�����z���������������������y�����:1k��?���]��km�s+m������������������������O@�Փ�]��� w�i��	�s�b���:�<���u�a~EPO�i��zF�׮����3_���������������������y��i�2�LS��>����\_��}�b�܃�<<<z   <<<<<<<<<<<<<<<<<<�nx/P�|]=M�ޭ���ϝ?��<�<g�؎(W�������Rs�D�+<<<<<<<<<<<<<<<<<<<<<�wg6�?T_��+�:�e{w�5�G{��F�]e:�I�^�;:����γ��%�����������������������|��P�fH��>:�㮾ª�n_�u�)��\7�3<'���x~�tȴ��k}7��������������������������uz�}b�Џ�X�<�ךx�����������������������<�sҟΌ�ʓ���Ks?����ws�s������������������������@���t��Ҟ7����'��%	#+�zޙ;���'xxxxxxxxxxxxxxxxxxxxx>�sR�'���}�I��k=�󱜮���;�������������������������3;�#�#=�N��DD�ZO�����<<<<<<<<<<<<<<<<<<<<<����w؝ݳ֩u���Y�)�����<<<<<<<<<<<<<<<<<<<<<��u|a~2��䎬O=�������w����_�yxxxxxxxxxxxxxxxxxxxx�9�w�<�3Y�.�ˈ��L��頿���<<<<<<<<<<<<<<<<<<<<<��^���1�uTbJ�k����uz���_�yxxxxxxxxxxxxxxxxxxxx���G:m�Δ����igt�H���3a�k*��������������������������d�4�Ԧ�:�>'q]d�e�u7�yxxxxxxxxxxxxxxxxxxxx>�s�-���N��wz��LXu�ְ����w�ֽs�x�}B�\t�tJ'm:�����ȇ��w�yxxxxxxxxxxxxxxxxxxxx��9S�'���#ө2�VLuĽ������������������������y��O�g���)�����l`��)z   �+��e��3<�k �ǭ;�c���h�e`���$O���6�����������������������3�$}��[�l闣�9`1��^��_\���k<<<<<<<<<<<<<<<<<<<<<�MV�0v@I���y�����w��:N�����������������������?�nf���ө�i=�������p����/Hdu7�yxxxxxxxxxxxxxxxxxxxx�9i]O�Nɨ�ܟ�����1�Y_#�����>B����������������������='��]Ϛ�^G�P�����w�}M��yxxxxxxxxxxxxxxxxxxxx��9Ʉβ���}����i�)ҏV��z�e}���N��[��w-�F������	�.������������������������8�}��ݠ���qd��n���n����/�>^����1���D2����w#|�z!�3<g��tw���o��z9������f�yxxxxxxxxxxxxxxxxxxxx��9���tsߵ���_l�g�'1$�{!�3<'	�_��9�N�u�dy�2��6y�Ɣ�<<<<<<<<<<<<<<<<<<<<<�U��9z٪�-��w�u�aOٙ型wY$<<<<<<<<<<<<<<<<<<<<<��\u�Lk/qw����;m�OE��/�Cl4�3<�h@ߝ�5�}W���Ǫ>w��κ���M�����EWp�]=�}���;��/2�<<<<<<<<<<<<<<<<<<<<<�����MY��߬�$�̇��_��gx�����r���~����ޙG�6���O�����g&���������������������|��H��8����;�㮾NKL�����u�"z   �G{N��Wu&��m�����ߎ�rw�5ϧ{N�^�z��>-�/���7}���{w�yxxxxxxxxxxxxxxxxxxxx��9�)~s�C�n��V{ci����������������������<�sz�z��5w���~�����6��6������������������������'�����.qW�b�;�����9T1��|��������������������������:Ӱ?�"����ÿS=#�kW}��������������������������<�s�4��n��_V��W�n����>i1{�An�xN7�(U���&wW�Vz�E���IK�������������������������AlG��z���U_�V���"��xλ3����h�i�ײ�;�����������������������=�e#��2��$X�����uz��F��fxxxxxxxxxxxxxxxxxxxxx>�sR(E3��I��qW_a�k�/���{�������������������������sWk<?�:d������������������������������y��|g�:=�>�_�Gw�u�kM�SBxxxxxxxxxxxxxxxxxxxxx��9�OgFz�I���v���ƻ�����������������������y�������0@��W�������������u2P���#	w"�3��u�D֝��ad�Z�=���9�ϯ{N�I�ζ�}�ρꮵY��,�+v@�?G�����������������������srbws$ � 5�s��,�B�At���_�yxxxxxxxxxxxxxxxxxxxx�����;v7F��u�zf��,�,�|���<<<<<<<<<<<<<<<<<<<<<wx�:�0�2���<�=�������;�D�k�5��ӟS�1�䁤�z  �o+Bz�ެ��$�o�{q�;<��Yw��:*1K�m����u�����Bk�;<Љ��:S֫:�7ȯ���%#���1e�k*�����������������������齻$Ax�������I\�~[h�A;�O{����N�t_�l�/SVݠ5�=���S�u�9���<!q.�a:K�m:��]��������Z�����������������������9�bOb��G�����j�#�w���
�yxxxxxxxxxxxxxxxxxxxx�����,<d��������ϖ��`��^�����������������������+�^�=n��C�$;�Y.��0�G��:`���������������������������&M�(��[��(uXLXޏ��W�V�������������������������Y�����(�!�왑�����z׋��yxxxxxxxxxxxxxxxxxxxx.���s�|�v�	�g�Iгt��]n��^�TVw����������������������s��$��E�$����$��.����d}��~��#yxxxxxxxxxxxxxxxxxxxx~��*W%?��\�    IEND�B`�xsr java.util.Random62�4K�
S Z haveNextNextGaussianD nextNextGaussianJ seedxp           ���~E�xsr mobs.Player�f�;�['� I carryWeightI dxI dyI expI heightI maxExpZ movingI nI widthI xI yL armorEquippedt Litems/Armor;L 	inventoryt Ljava/util/ArrayList;L nameq ~ L skillsq ~�L statsq ~�L t1t Ljavax/swing/Timer;xq ~�                             w    x                                   `    psr java.util.ArrayListx����a� I sizexp    w    xt mesq ~�    w    xsq ~�    w    xsr javax.swing.Timer��	�8�� Z coalesceI delayI initialDelayZ repeatsL actionCommandq ~ L listenerListq ~ xp   
   
psq ~ ;pxz        b�PNG

   IHDR           szz�  )IDATx���O�w�YBF�2Ra	Lel��^J�b[�-�ӈEZ�j)�R(�8���V!�����r�`1s�K�Nd�v����2�8�-�٫�wO��?`�!Y���7������s~�9OH���?���Y<]~�_�������X^~���%<~����u<$���+��_�$����w�'������U�x����U\�:L~&�.F��1==�� ���1����(&&��>ff����<6�6���	�f����By�2�T��_\��on���׋ߞ�`�E���w�|�2M�k��O����w�Ne����aܺu>���������2�9��{�����B��y�ػ!HK�Å�N�'� v���L!$�ݐ��������KQ{L�#� .�}�}�y�1����9LNMb�ㆹٌZ}�ǤtU�p:��s���-�!o/=;�hM�F_�%�r��#l6p�\z���جm()U!99��&<Z}*�
V�L&LfSz�2Y@�<��N�a� :�j�4-���
+����P|�o�� m�t�4q�L���$��z3(��0@�R��e*r� ϑ����XS]4��`4T�T_���x$$���n���[p��i�@������e�4�ZS	���CTT$�Q�))o����Ɩ\��ِ���������R��rt�7�J{��_��l�=,ҫ[
���@�wjE�xX�>h�֠����� ��õ�XCQ:\����=�e�E������ @�Q�L��X�y\P�c%��ُ޳֭��m|��4[daa.8p����C��#��&������֒�
��΀�a�(̇�\�Z���2�������Ja"��n��L�ok#�C�z�����B��H�J��U:��8ⶩ\:��Qz����=J�Pdg>&}'�g	��N21�K/�reY���ڞ�<y.�D�Dý<+U�@Lz   ����s�i�">���<�ތ�&������tv���D@_U����'m�h4ב��}�L�+!���bbb��N(�fo��o���zu3 ZflE    IEND�B`�  h�PNG

   IHDR           szz�  /IDATx�ݗ�OSwǝs	Q,���J[�����aC\(
F�[jK�ʓ�YV�<��`���A�o&٠����mऄ	0�@�W��G��/��l��M�9��9�s������=[ucqa�[x���}_|����M������W�;fa ��7��ӧn,/=���������˗��j_������y,���Á�ma��FMMF��K}���0==�É��f���6�++p�f1>>F=��D�5��/���=�x��
O�����=����R�j)�l��|�p
c$ӹ�9<z�FGG1K��u�`bbE�
e %z=-��I������Vk::lhmkE�8��Q0��R �lni�X,��������@�DRR�=v��y��N?x����"8���xP[�����M�G��y6�2 ��x��d�Ud��� n\J�A���vle0�0������i.+���RTWW�ˍ��G�^��
ȕ
0�LjG��J��� p��pP\l����ɻ⋔���U�
�����C*���f�Ώ$���لxyy�4}�g�R����@�G��s�+�!4,�ŉ!
:��5ǐ�(Ftt$.H��l�"G�1��T0����{l6�T���{�{0���G����@��8��`)����M�
�����
�P�;mֽh�Z `�x��PK�	�ӓq�TB)��;�����f3:m�{��(�o�W�ǋ�N��k�:h�0�5ȑf�V {׷;��U{ ǝl�A��./)��4#�~���w��{{|4�Z5MhQ}��\�2��r���J�I	q��rA����?����Ib����.�S��aE}M)��|$B0I&�����|�� �I�'�z   ���m�u���W ���c`�8r������� ����P�A�4z��&\�H�6+|��{`����0��-���x���Q�=���ݝ̌�g��8-���s?�1�S���>�6Y�ȋ�9�YA�H�UU]A&�*��T�Cػ�10`�`�G,����2���z�r�d� =-u����7�?ܰޮ=    IEND�B`�  ��PNG

   IHDR           szz�  OIDATx�ݗ�O�u�'�A|�A�2��
�
�R+
�����{c\Z�[[(��&E.�[e��0¢5�{��$�ư��FA1{��|j�>4ѿ��Dϛ_��/9��|�y��=��W��/�X�|�?ކ���4���5l?~����w�������&$�[C߃���_q��Cl�6�r������]A:���V�����8�N���K@�`6����䫰xm�_,c���v;�5�Z_���l�����5�֊_߼�W��j�b��:��}߮��YH$�Gɓ��n���>:p��W������>]��e��P�"V���T3��������C������v� ��l(�ŉ�t�Ԩ_Cjj*�A8q���S`�"--#�p8�ä��j�^�mr�~�g�P�bvn�,&T*%�E�V�h�~�{z0}qW�+P[��@?�:T�Vdd)i �͵���4j�0!�����H>��B�p�y�TD�b�H�0;�	Avv6��R�!�"66VOZp�Q�W��*�J�ti4�*ĲX���@\\\�ĨY@
@C�\n,�����`��FNV��<���h�m��_�KKK�%%�p&��\y���$Ԩ(� ^�SG,Ú)�����6���d��:u�填�	%�8r�0"#Xe�65�� ��e����'��E���$.4�rȤB"�ϸ�&�12Է� ���'*. &��v|���2)��h�(Q,<����8��ݎ���z   �W�M}�T_��ƺJ�y�`3|q� ߣ����1	��2��)��tĔꣽU��bj���_	a�9��r������<���o֐�.�h��(;��.��3��#22
�f³N��.�F}#t-5�J
���|��������������۫��O�X����N�$'�A�N���Bazzz�JZ+V�d�5j%��x��K���E8���_H��JC[=
��;�짥�����������������=��)�����2~nmnBUe9��r�U�d2�X,=0u�0��J=nS�(WɈFc$��E��J٥�i���̯�����@�&]b=    IEND�B`�  h�PNG

   IHDR           szz�  /IDATx�ݗ�OSg�YH`�%�E+�rm!��PZ�[+�J�n�p)Rz���U�6E[l�:��e\$����K�y�2p�An��&�-F30�H�_�K�=����&���>��/��j<��nݸ����)Ϗ;�����>]���,�/a��u����I��8���X^y�ǏW0?��ŅE<\ZB�P�:q������^<���e����/����t���%_�7ob��4�������~~�>��O��,Y���v��o��O33����p8033��w���.�^"�bi����~qw�����8&����+&&&py��&�71�F�����s.��͆��n8۝�$#%%�l,�ǟvtvB|H����a�Ex�^ĳ�!�amm!`�7��Ӿ�����2�$�2g?�Y ���[h �Ԋ�>x�����цv~���B ���רW�i��zlv��(�h�͆�@
�F���U��frd�A�d�4�BX�.TWW�d2@#!�			08���F�^T���l�A*݌���`0S.Ws �Z��^j<�H��r��0�S(�-��L�>�X,�^�#cCv���'��F��>ȅ<��J9�� ~~~�������,�z   ���6"�g��H�K�	-�C�5k!/-�������������Y��ܚ��㢱� 5?�"��-�7�:\���8eiZ3"�����|�2TF3q���T>����o�)�p��x{�R���Vp�I[��Z��Ӑ��,&B�~s�	Պ�?ʸh2M(�dl>��L�N[	�(�>��((�C.�BBB�p\K
 ��cd�M�F�A*}�����8C)�։ ��y���s��v���P74�2df��No@{h� :^#�R��t�rz��AW�iXj�E��
DPP��`�J%7~���[㫄Q����&pR����E�%T����!�����Q ��fM���s�~��-ũN"'G�$�lFF�18Ї�v;.�J�`��52��!n��jQ��,$���%�̯��>��/:D ?��    IEND�B`�  Z�PNG

   IHDR           szz�  !IDATx�ݗ�O�Uǉ��R�Q7�t�ɥ0Ve\lR#B[�K�h�:z���q�BKmi�:�u1�Έ��̙����ˆ���2�E�_�/��b�$'��$������9���Z���7�������}��/����+<|����e,,����O�vn�`�Z���_q��f��q��]<z�3&?��> �w�`��%ܿ�fff�����''a�Z���J/ĕ�3�ɩ)ܜ�����`��~O�� ��0��趛1���9}���r`~~ӷ�������W�>�{��d×���xp�����5�32B/��F�����Mp��`���崣�ց�H8� ��uİYYY�#�<�^x�i)����H%������߇��\`��j���Z��@W[�6�56���t�
a�耽�So���0���&1t\�D��I��R+a���B�EB4}�����(��d��[ �U@��F�&@xx8} *���i8Z.�N�z   �SO>qI��*��삯�/����nj�HON�b��}8��M�\n�6HHR
�_������-�;C��|$p�Q�W@&-EM�TU���f�v���k�����#�b�;33RQoP��]m�ǥ����7�����8kn^{��gmع#�Z����V=�(/FY�}6Ps���\�C�a��rxi~fv��P\4�c�LIđb�
�iӆ�չU9�4կ-�������2����jH� 6t+8�,<��B� �H�d2��''�}����']�D�G=��a:"~�I�͎��Q^I�"6KY�ǱO]8���(+��&3���Z???�����Cm��n.����ټT�Ehh�!� ��b[���th�W!��C
�	#��K�����H�a=&&��b���Ctt$rrxrZ.\�CP��m�S���֬�EEEU�ʉ ) ���k���Z%�:�Cn@/Q�Rr��UB x�L�=.�v{;��ۼnO��!7�������0�����(�d<�����    IEND�B`�  E�PNG

   IHDR           szz�  IDATx�ݗ�O\U��Ј$ZR�C)+P��R-�!¥�\
��0�� e
J
B����ڦ1B4�Z�����E+�`��j��<3^����$������o��>�v�����W�?`Ux67��'O�1������K���ۇܞ��66�x��GSS;1|�"�w����mfg����[[[�������W�7��9�ss,--q���;�477<U��׹v��ϸ�����:�~|į�<f��
�O���+��:MB��k,޽���2��_��p��#o��PSWǻ�]Ƙ��Ofcb�fff����!Ð� u�:��9PP�����^��YGsS�G}������0�B��j*#�;qqqt�ڍ�H.2@Q��%<<&����c6�u2�3���h4�hH�<v��99�x
)hFW��z   ��E�B\ ���z;	�j5�J%~Ύ��j���� �Kpp0Z�V<������}��塪P����RTe
J�[��₣��x ��D��RX���\����def���E����R�͟f���Q �\������MTd$1{�!)1���S��99bc#a�-�8.��F����Y�y^�d�*NS^��Tj�L���V��4l?����I����DH�K�T����Fey!��b��,�H$��n�՞�~��k���J��ue1j?O�U%d�J���Y�ZrD �]����V/�k�2�}�$T(�Ѩ�(��"��P���J�k9ǽ9��l/�����?�����h|OMN���'��\��{HII"#=�fm���d��}[|���|077����h�V�M��'�v8���ar3S�D���c�W[�5p�Q�B�MFj"��899��677���>8���/�ML\J0���T������#�<�� ���&��@O���� �F"ٙK驌����������?3��E��(';8@ȹ웿?=�(�'//����]ho����D���$/T����Q-��0����c#������[�(�C�~ۑ=�ӣ炾���]޹�����yM:q~5�    IEND�B`�  J�PNG

   IHDR           szz�  IDATx�ݗ�K[W��i�b�S|��K�I�,�h��Tg�5�j�MbMڨ1i�Ƹ$v���N�01��QcײY��.S�p���V�lc?̦2�/�/�A��8p����~��<��܀�����x��߮`ks��;��}��?���ί��s?��{�W����Gs119��/f����������nܼq0 �����|��~���+^�n�n�*~����+x�l���a���ona��<x� n��^�_�Ws_⻕Ul��	�׋��u,����yLLN��h��{܍{S����H��1����<�S����J�5�XoA*-����L&8��P)N"�ǅL.���z   �Ꮗ�����<~��D��������h4�`S���c���[���fG�㷿N"nQ+��X���Ơ?&��	��コ���Dzz�u�Ж�aG�Z�r���連�cb���!��X'*J�u�d4�iD�R	fdZ5J��'��dzɤ@�Q���
m� 28�:����q��		|�ǆ���j!����*F0NVW��M��&�d���A� �ǅ��J�lТIu��c�oVè� 6�6;�������� Ǌ�&��D��V8��8�o�Ť��<0 ���r���]~���#��I�r��Sy���&0�T.�8122B.�s,�x,��&t��h�¨S�Ht�_`�~N�.�ſX�/����h�_���L/�+q�g���� *.
�PY)Ef��w����.T)贙0���T
��HH�'9�#QF:BCC�_#���a��d/v���w���@�_�ZN�#�hHHH9-����S��0�ף�r�� ��-e��H^6b���k�P�j������.�ڴ��^ **��b6� ��jP��cG��7��"���銋� �0o'�_j�6��� EEZ���ᓑ����M����]�D
�юW�.�����ߝ��
�FD׬�Ym#� ��k�}�L����_� �6����    IEND�B`�  a�PNG

   IHDR           szz�  (IDATx��]L�UƉ7b�e�����ʆ����Á�Q�G;@�R��5
-�h;�b'�b�!&Z4��0�M�0vat����7>�5�{�����&�����;O���_��bmnn���2�l�я?aw��M�n��oc���_������G��������ffgpX�j	���������� &��g����˅l�����a���E���͍(�v����ְN�w�v`���pg�das�9;�_�օn��1�Á�[��X�ڷkz   XZ^���y���Q�%�B�^LLN`a��.����2fgg1=3�y� ֮n��� 5E�F�ju,��LF4��2jL��@(B~R���Z��riii�2��VC-��m9:�022��I��
����!i���z����MЇs����uJL���%I ���@-� *�
�G`4� ��e���	�zT�"??"��e ٧E�ՂcP�� �I ���r9�����:e%Ȗ�@��B*��I���"��f� O��1�{�� ��M�H�E��˅��"
���A�Ét�:�N�2Y�45gQ�*F'+ ��
hkU�����y
��� ��q�%E���AB<��*�G�:t�
��3A���11����Q�C�v)�w+�P�T9o�!�7h*����Aw����;���x���Ҫ�q)���I�z$�)t��$���9���0>�k4�K�EV|8̆�)��\���N Al\�7x�@&���/�L��F���!�e♙x��V8n��}�i^n6�j���j��,u������iș�C�`���T��6�FGQ&/D���}�����ϕ싒��R҆xd��� E���C�>���NDF�!Y�䞡4G�:r$"����,-B���7D�����b�� �����\6k🽄cq�!H�8PY��E[���
�����0hk5�d���M�dDӢ�I�� d�w:03=���U����S������-.���rVX!!+�>�Lߌ��t�Ʌ��������7��>@���    IEND�B`�  Z�PNG

   IHDR           szz�  !IDATx��L�u���` [qx p��L��CA0�#䀃C���8~(�%?dNE�l@�ďLKS�F4J�sKm���s�z��[��s[[���w���}�>���y�y,�/ֵ��鱱qfo���{<}�����t�>=�������$w����o34�o��w{fbz   b�˗����<y����.� ������;��0??���(�_���}��3Qś�\�gf昛�:�#����/���]\�s�Kܘ�嫩)n��d��<��_p��:::�8`����Ӽ����/���ə�3p��s������+��B�)�Xc�`a�Щ	�I��U\�*C-��ꈌ�D�
���� 66�'�����</�z7g���a�0x��ǎ�jj�`���\qJ�z4�7���͛�Y��Z#�%���Q��P�)�(������d���S^QNe���U+P�f����0��[E�br��e/8��j(�W���ԟM�6��+t��#	Ev�w����yz{s2X���{{;z;������b�a!!�d2�w ~{�ի��}�����踘��-�P����K���P�x��=\Q)3(�߃��/K�qrZ"�QUU�`q � `kk�~���<����Ъs��H$�<<$<�p!��t˺p��O)Ӫ͇zz.�D��4�OXsQd�"qv�o����-�'.n�eƆ�(u7��с���]����������\wss��Ǜ�0)����h;f���|�7WA�e1R?_�c�̳��Z.�t82!+�J�� RRv�v��=~�^������
��KJ�cWr<�!��	H����������pɞN��N����t�2vR^Z���S$�o�����]��߂�Z"����� ?��Qd��TKhhq�1��&L��!4d=��˨�,�S�靃�\�'cا"::�ۈ�`V��~���q�!�W�̖����RG�NCLtԳnO�5r2b�uF�/+�l�)Z��	���d,�@ii!�o��|���9������V�j�y��'&&�FsK%�4��Y �KM���P�    IEND�B`�  N�PNG

   IHDR           szz�  IDATx��YL�W��h�
e�Uf�Zz�Z��BՉ�2,3:0P����,�H) #�Т����T6��-�Z�^��HIz   �Pӄ+{��w.4�l�?I�~����/���=�{�������ҥ�џG���^����ۃ��\�����_������SLM�����F�% G�}���,���df�!�����n� ���19>���[�������C�������{Q��9v�fo_��Ì	
���2���s\��5M�5��B]]W���y��C<��ad���9u��� �G��ɵ�ktt����FgW'�����ζ�����D�Z�����G��s��H�s�Mtt�� �`6�Q�IRF*'1:�$�:t:��� �v��^��D�T*�>�^�w�?Ԩ)6�`�Y)�,����l��^��C8�:L��g�(�g���bJ,
M�ą)�ZKٿ�N�ď��l��0U}߸$�)���=,XH�р�d/��$lڴ���d� ��R�%��c0�
���s��eRV��f��Ex{y�}�9P�G52����mlyg	�^hw�@�5�LJ�B������$qT���F ����r2)��L�!�|�N"##���T���ϏO�����[����ܚ7�(+�&j9�E�b)�G���yc��Kp_�"V�<�	��ùiH��}&#������g�(���ۋ�E>��/@���/�O�{8^�sn�訥��7��Ē���@�K^(����	\�[�h����p�8���n>j������E���B��_aED1�˘G�m��/����d���˰�l$��'y�ۂ6���g	=<<�1̣���VE�dKB(w�mĿ+Xq3a�Vٹq��� ���P"��cEh���|� S�9�cMu�ǯfg��5=a�j-��D"����U�"��O���l�+-�ClؐDԲ��g��ų��W.g��8&:�.K��Ȅf��� �'�����#�X̜?w����4a�;�-�ص;��Zp���
��ŋ����f+����D�L�.�˜֔J�����5=J���2m    IEND�B`�  N�PNG

   IHDR           szz�  z   IDATx���kLSgp�m��eRN)���e��@,�2��@i��b/���R���B1�8.��^���	��2p&,n2�2A�H�0�a�lf�D��^�A��Kz�,ٛ���/��w��y����:�<�ǃ������u��m�6� ���2VVV���O�,���?�����t`}}kk�cu�W,<]�ڋ��=���!,/�`yi	����=������	�^�3��g�M}7�7G�����ssX�e�&S�U����޻�o�qwb}��`�c��O���qW�^���f�͑���̌3���p�;p����>L/ ���	�������f���%�=�ٍ��Dz�R���x����+��;-:���TT��`lѡ���8x0��PVl�k8%��ώ�P��a�쀩݌��Lw��b0�k�<?4���W�����Г�H{?Z��y��(�T
zŅ˃�d�k�m� �R������<(
������Ł�"#H�

�oyx�����zH8l0�L�X��`i7���A&�Aݨ�n�wQ]Yee)�	v"���A�����ijq���D���yf""���͂�?L_|n��������'�tJ���h�J4��@ CQ���A`1(�件
sS2i�sR� �LL@�a<j�JPQ&EQx���,x�s~��3��1z^�trr��:��+8�������ΰXLgR� ��u-�Ԫ}�`�>��:ihEX ���������E����a"[u�R�TV�nU�ɕП"����bq87�%������\T�?%� o���B��%����o�(/�@��A�3`4����A����㎹\�6�m�V��`Dא�uU2��Ga�ԇ<q6�s��M�J^š���1�4�U��ay�j?fm���t�#�J�� ����{�Þ�����$hnR�Vu�5�|�J�q��M������7�:�	Z4�$%'��LJ�.�ؤiؼt�,�6�s��#z   ����(�w�����f��=��r��`;�O���    IEND�B`�  4�PNG

   IHDR           szz�  �IDATx�՗[LTW�m_����\a@��X��)���2�6(� r+3C��(3�Mn���P"�M�hMJS�)�(/%�H�X,�4mUlI_4��qI�8g��NN�����^�:�l����̴i�����f��r�V���/�a}m�_~����"�����	v�����O7���#n��1wk�ǏVY}��> �==�Y^amm�籴���l����/�&&'�X���e��O�<��7�_����zq�0���Ս�7Y^��7����066���mff�g`pP\��zW�\���q��gZ�Y�q��kSLM}���Qq�ԅD�������t�^�9�h���Z�q
�� 5�夤�����;),( e2�:��g�0U�m�����A�J%Lp0����h>z�ҲRq�չԿ�LәfZ�Z�7�J����w��(���*.@mE1MiJ��j�OT���\OS�?�oĠѨ��;�ެI��X��P[C��u�:*��P��E�ӑ���(*���H���hy��(*Ҡ����T¶m[���iS!!
����-e��%:U.^^;�����Dzz�8��Ą8�:nnnd�#����E�"��w<==��n
�9@|�>���Hz3��S�i~;��UZ��E(�����] ��舡��9?{m��Tc]4<<�����8*���=��988��"A*�NFF�mnL|���>����|}�*�ޞB�";�^.N�������YbmT�������1&''����Qk4�L=�Z�!��	gg�__|}�	�y�!�-@c�)~�|��(ذ�3�m�D�F�dr�!X(���J$��<�����DD�臥�����C� �\KO����#,is88J/�'�n�)SPdb���P�Y���FE���Ņ��H�Y\�l�2����J��Ňx��������|7�##��HC���Ǣ�
��z   6wPUY�	`2T`��<kF��n�6[�L�W�} �+�����قJU�dwqCM��GG��R�P��dA*��������.�NE6,    IEND�B`�  U�PNG

   IHDR           szz�  IDATx�՗�OSg���0�r�Q�rHm]�b���Ei��P`\�B�Q��":�\��2�l�6��@�K�l�l�q�)ˆ��8ْ���N�@��4�I��%���>��w۶�վ���i�w��n�|ٜ�Q�W~�Ɠ��_�����N�u���[��W,..a��e��y�J�ҏt��ݸ�z��}�M[__��lµk��Gazf��V�>�add[��G��p�a�d&`��s������s�X,�������.��d�\���o>�x7fg���
�}��;07�((0HhkV�?6W޵`hx�WaC��g[���R�4��T5�r9�����>�6����dp8���s:���d�]�����}Е�1j��T�߬"@UYb��c�Ytuwa�j��]��Y,�28�\���4Xu���`h5��;��|�%�A���(�r$�oY�Ң"��4��L�Z��"��b0�Lr!�Gy��W@��Ǯ�@'"PJ�?/%~~x{{�������B	*++�#�׉���"**�������@h5jd�v��e�!ĄL�t��` :&	{���������Dس����0y��СQY	:-T*50""^^^�\&q/�������Z4%y/������E����|�����N��q/��g��(�t-�U}���h�֡H"D�����Exy����:�����w\�f�3�7��C3!+.�e
v���0(�%��4��Фӹ@$Q�m�O:���$l#�C�Tmc��j����nvv��$����F�%�$'���RH�!|��������czʊW3Y[�
�og:��C-�~�W�z   (7���lH�Ѥ�A��'N��Oi\|"�">n7xy��Y�b1!9) B^^�(b8}� :*�!�s��"�9x��z�Պ-�
�SO��X,}0�va�6�%h�x���g �$		�ټ���F{���Ty��h��||��F��F��(�ߜ0))q��<e���7L�Z͉    IEND�B`�  b�PNG

   IHDR           szz�  )IDATx�՗�O�UƉ:�IJ����hK�J�Z��p���2���Z�ߦЕ���V���\�E��l�)�-#�n	�����˂��Dc0�l���?��~����$����}��s���ך����ￛ���*f���yV|q�o���{X^�������*<"~���6�ZYy�����������l��!�lm6�!�[�[������_X_[��a���s̻0:6��o`||�W�`��M�?z���)�|6�, q��goa��M�]X�ș3���q��-,,�a����
��o��:5�ɫ������˗\NL_����|�Е����Ƙ����Ԅ6�==N�����J�:Uc u����n���"N$�?�� n b�� ��0��0�[�i1qۻ�0l�Eo_/~q�b���
gxJ�%P(d���K(a��pv�cph߶�Y�';Ob���A���07�v��TY�j�ٕ���H�R�fe���E^^^/2E%���Ʀ� �Ɉ�b522�`����EqP��C��B$A"�@�U#59	>>>ص�%|~�'����:��BJ�/(!B!
�����|���Ɍ�:3������|
y*�:�E
��Xr ��P�t:f 4j
���O���a�)G��}�V��u�G�`�X~|�B||<�c$Kn�vn�)�R�N&!'��Q���k�L4v�f��BC�x��}-��0~~�oq]���y���Q�G{s��W_V��&��%�d ����������4:��/R��D�-@ �_�����C"z   @8�s��6񴴔��$�g�����I�~jU>��i��)���CɈ��Erb����ͽ{�u��PNk��4h-��B�І�j�HwD�"<c$?0��Bn��(8�-f4֙P@b�r(�����G��`� _���Ϗ�2}1Nu�� ��BIJ����e�P��rv���Q��B�.(` 779�� ?_������g�t�N8�:v��J�Po�@ֻ����!4�4�sr2����ao��g �_�r=y��@wL�A�y����Br����    IEND�B`�  V�PNG

   IHDR           szz�  IDATx��]L�W��	Y��YJ--e�m)T��Rk7�W`�!-mWE�(�:��Mbe0AƇa`�	\�^Mq
��ɔL㰛ܕ��w��KxI��$Or�{.���?�s�y�������\���;w��O�k*>��n߾���_q��������ϯ�����Ǐ�៨�my�Va��Ct�t��t6�/����p��^�=\[X@{G;�����)��O`rb�f��>nݼ��+�1:�	� ����Ə?\���ƃ����"����^��&�����8�ù��03=����1C�������,f#�.��� ��h�p:[�����jCJ�|� �҂%ZZ�N�d2��pXE�!𐖖�I7���
�jo�{�La�Ŋ6��񠫲&#J�-�4)�Ѧڋ�����AO��r�Q\��[Qd�+��l�B�����X�HGC��^�Co��@�ӡ�^>�O��T��b�r9֭{�>��v�+11������*��tP*���?:;��h(+-DR�v�:�N�p&��p�d�!����ذ!�=
z\HH����LV������z=*�2 ""Q�\p�h4��hn���l6擓���KPEď�a�(BHH���`���X,�V�Ԭ*@���'\.�Z�4Q����pԽ���B>O��z   ���jQk,^^U�j�����O�eP �l�f����9��ӥ��4eg|�j�MΙ�7��fHK(�m@��!/�`�� jn�)v����Ϭn��5�<�ɃP�9�{9�H9���|��&��ܟ��(.=U�93�m|����
նrI�h�+-	[X,J488�ҦM/^��dݫ���RiB�݂#5&R�D<�\Ѣ�y��*!,l#8�,TYJ`5�@���}JhI2�0p�	[�`26�ϷW;axi��8P[U	9	�FG=<��R�mAG{+�^c}*X[[E�crs��hhnn@w�q�t��b�4�5��Q__���.����yq�+l6����YGS=�HII�����/�_�1c���    IEND�B`�     F�PNG

   IHDR           szz�  IDATx��[L�gǽ٥a�Nt#h�3Hq"gaTE�R�s�@�C[hAZ��LQ��eq�4��c�c���-��m�������n����I����������?۶��5262�����_}��◌���޲˿[���o�q�;����|>;���"��W�r�� ���o�|�Γ'����3�=��WV���@���r�3==�ڣ����_���͋�/�p �V#.ĸ�33����q��K_���hӒ��y��Nq����)����Yo�drj���Ç?���$�}��(�ׇo�3�r12:�ݏ�⚘�������Tiko��a�A\8kd����BW���N:?��f#[Ntt�l�T��0a����7`l=K����s�GO��<��V� 4եh��k5(O�PW_O���j���FKj
����n�q����24�
�B���i����YS���OOO�R)2��[._h���HS�^ hD]������*��z
��U弗�L^��$���,�*RV�;��`�Vk�L]=F��N�\.�XR"���U�PV�����{��ߒ�
sS�J%E�S�
݆܏��ޏ,=�I���=������z   ��)x,��ň����	G���%)d�C�Ԩ��D@@���}��XÑ�qX-M� �HKM&NKLT('d�ߺJ``�8����o�b�Ʃ�47�8EDD8�a� ((H���cVy<!p�x&�)�������.�w��}�v����������n��T��9x��o��l�����;��l301:@�2�Yo�ҽ0>N�y�]m�Ǹ��~vKt�?��PU���Ĺ#����htD8������A���p��u�Ǖ+�����V���9IffQQ�$M�@�G����9�§*+A!�݌�RE>�3�a�7l�������~ǧ¶̂��r�x�ߟ�r%�����J����T��!+3���D���`�Y��5 ��J$B�J%���V�����wǥNL����xk�α�� !�b����*��FͶ��U�Hc��*"�    IEND�B`�  m�PNG

   IHDR           szz�  4IDATx���O�g��ESn$�F(����8L@�e7d� �,2��� �0�2�`p� T��i,%5��$6�E5z�Ҥ�Ջb���O��Ĥ'9y/���w����Ƹ}��ϷO�r�!S_ܣ���iÊ?��)K��34�9/~}���Q�ls�-�OD/�����f�oVVVX�s��[��7���?���iDh��3>>������`u��~ͫ���AEe���n��{d�K?�ĳg?������4V�U\ ۜ���G< ��gǅ�_���?�/@II���.119���A�S�����x���P���;e�D����|�n��־K�7wg=�VNǆ�i�nj�O��k{3��k��&�z��78w��vs;ƆzZZ��(W�S���JUN�Z����ZM��,�-͘�B�'D*�n��E#�u�)�)�Ҡ�ʦF[�N���e3M
955j�b"qqq��Ǉ��4�� z�Z-X�mh�(*-#7/�ʪ*4��NfQZ|�����3����b�?�^�JY�z   �=:C+��V::{8�Ւ�_@j\,�3��g 3vFC-�����D]m��lR����D&c�������ۛ�c)hkTtZxxx���;q�����T4ԪٷO�ɬ����ř<��^���ř]]�zQ��^�($*z?1B�/���6�ƭ	1N C���GRI?v���"�B��H� �IIIN$2"www�h�AkN��bb���K�?9)^��-8;�/�-���!�LT�Nrゑ�{���$~���w�2y�*�P�T�o9�qk����O�d���o`��i��0����F���2ܷ�ӥ�\�~��� ��/_.���(R�і��|�+���1̠���r���	�ͩ)W;/�A��;9m�J���݁������,,| ����s���rrrhh�100�d����룷}�6�������T
E&Je�/랡R��vV��%J��]v킫�������^n[8���������,F��D��pOt=�yB��#d)>c|�&z}���Aoo�ƈ22RFtL2��݃�'�8::ns�?ޖ��cx�E�G    IEND�B`�  T�PNG

   IHDR           szz�  IDATx���O�g�I��«yA���EX�M���(����`�Sa���
�F9ԁR2A7ġ8�����酧���d7K&s��y�>{�����$&�%o���}����}����yU������#NC�Mm�����=`e�����/���m�+6 �֞�����<[����v���r!z�{�_�ĝ;�y��/_����u���8���**���$׮-r�7_��|+�����<��ss���������W7�X�q���\�]LOO���*��d�x ������N�\\d��U�\a��߯�r��}ܷ�tuw�0;;���i3c�gfq:r�a��Y&&'أ%,$���� �Ǉ��a��a�h����sG����B��:�v���9QL��0�uu|��NUu��V��؄�z   ��Rڵy��
��^p��))ȧ����ړT�j6@<
�I�ӣ���HXr�*�j��Sd|��a{��VZM�TV�R���P����J�!tǉܽCQM�:����kI���in<EWO?�a���M&�[Ա1T�N`�Ɠ������\��3a4�D��C̾w�E�O�"���$������,���V$Ɉ��y��Q��&r >���2�"d����+/fD�+$D.�D�������b1b�IH�#)� R_��F��X���!�!\������3�\T�	��Ųe��BwP�+v"^�*�i�������@�Ʈՙ�
ͥR	~~~��~�2��D�������wI�Mb���D%[�n��^p}��S���3�DG�D���T�/���?�&��Bw����GS�)�o^>�IW�e��f�5�d2&M{����Ӽ9
���<LOK��VG���ث�l�͊Z�b�4��R-̸���(2Ti/���P��qJ�����=3�ŹK�g�ܹ���
��Jy�{4G�w9�."#�8�'>.�cG��t,�`��Ԕd������WF����m~�ry����D�����oQQY�����&�T>Y�L�J�����՚�x�����>D��V*c<� ݴє����!�����տ�
V��`2&    IEND�B`�  M�PNG

   IHDR           szz�  IDATx���O�g����H���C(u�����B�Rr,H�Q@)�Ji+hP@�(4K䰁2:� ���9��D�d�b�̫e�����~$&�&��{����>��>NNo�&��]f�f���ol<���~`��3v~�������v��~( ������y�����vx�������������������^�����!�6D�}{�ťE��VY[_g��&ϟ���
���b��ŭ½{wY^Yd��}��2?�/67��z���2��x ��7G����35Ń��|��k�>�f}}�%�x F�����n�djz���F�z   7����2�%�=7,ħ�1�mt��h11w�0�L4�����a�Z�x u�R\X�^�L[�P[��È�QGO�����
�ju�( W����f���BSQ�V�L�������]���Ԉ"�2���Je?0��VC�z�F=U�5���45w��4�˩�,�Tt$y9�Z.���{��hJKh����Ս��
��K�����֓D݅J�K�IUDc5����s�=ah�G��Ap�?>�R$�((��!$PFFZ��K�5���^u� YJb��P*���� Q0��.C�E|���Ԃy'���⼈��Z���B����!&&
yl4Ǥ��H�����%Q Z������C���̌b �����0!�f�R�x���g���0p<$����ӕx�sT��/Q?%y�Q����ί�D�1��G䅻���;��nٯ=.�e��������p��um����h?��~����273���d���嘸���<�X��:�$55U�S�)k�*5�r����� z���[��z�V|���|rs�9���`�22����"9QAu�yl=��_����1aw���~90��d�O'�LI&1&�{����hJ�IS*�+�V�ZMff&q�X�	����v}������&�?�׍�#�(�;Ý�'��d2`��)//mo��𳨱D�� 5-Y�"��D������da�Ҙ��Ug�������z��/ &[GM��    IEND�B`�  J�PNG

   IHDR           szz�  IDATx���O�wǹZ¸X��0���9�S�"2&����3�؁���Bi����8�f��3F�lqK��d��]l��^��mb�'y�����=����m�����]�,tvv:U����,=~���}����i=|��l�w
 ����+/WX|y�g�����>Dom3q�����Y[[{��+�W_�r��yJJK�
0�fjz���o�q�&�޹������2W�]�f���������z   2=3����ܺy���'���12:*���P�����_�"�O2;������OO��ZZ[�0��Z�l���͘ `����W��q�]&h���7����1f���c�L�C�����)�� 99�V����&� J����(�j4T����jj�����܆y�6���`1գ�H'3S�J����F�@-mm���VO�*�ٵS���'c�i������r�j�(Tk9]ZNiYC��Ah�
8��$����l <<|c!��'�L��;-4��i4).֡��C�>E�2���ȚZ6>%�5%d�������"�E�-�'0@B�\Fm��!�E�z0�%2"�!�?F.��D_H\�v"�GW�KOW~~~� TWh���D���P/1�wLT?�q��v���+^7*t�K�)�,�رO�����R�?I	2$��;��'g�@4Zaa��"�/��l޼Y���OzZ�0�	����=D�����5�)G���7��q����zѪr1��/v�Yv�H(
s�]<˾�`~���	��O���{x���}=��O{�Z��r"#� ����g1��s��N���C�.���~��V���o�68D�������6;���１xJJ��Hu�XY;����]�wq�3�É	d�B�զkT+U!'����cF�g$'�S�׾y������J�"��	!����B����h��N�A���ٽ_�e�������ex����uuU�����p\\,�s44�o��F��kN���6�w�-�Es$9Q(P��\\�����|�`�H���    IEND�B`�  t�PNG

   IHDR           szz�  ;IDATx��[L�w�M��%&��L\6t�j��c'a 0Dm9� --�C[k)��8*$�
#�v �(��%[�S����8��L�6����ɮv7�X������{���{߶m��|���n���eF��li�w��Ž/��'x��&''���Z�[�Do�����z   ��g<y����<��1w>����"CC�7a4U����իK<}����u����n�{:;;�����
0=3�ܥ9>�urei��W�x��nݾ���<]���Y���zay�ׯ/�t:�3`��������5W�]cdtD< �R)���p:�q8�_\dt|�%a�0;礡�Q<���K�}-t��Bo_?ͭmt���������~<l���F�����r�=�X�1�LX�VtZLg���+Ш��9���lጶ�¢"�LFl56j�r�\\(�+�s(Pl4Wi�4���l���2�����]�P(�2��Hok���J�9��*TEgP��ח��てX�єx�'quuE.������\Ι���o�ꬕ���*���+y��OGSX�MGk5���u�n�T�Ay�8�aA���]��͕���A�Yo�#6�d�|2�w����p��h9a�!�)����H����ý������ ۷oǠS��$��q�.�'55�pB~ E�1�7���#�m���� �#7�4	��ϡ�'.&���X���n�v�I}�L���}�����R_���ӎ��P&���hR�}ij���PFb�;R��[��\\\����Tk�l/7���4�XL��-�eia>q��p��$\h!88X���ñcjz��ٹKLLL266��֟ߔ:~?��o9����j�g��c`l����0����顱��F˱�4ǒG��9���BoOJJ��o�_��T��������FvV:�����d�7�tQ��Y�n����LRR�8tH�/�����bg���s����dR�|���$#=��`���?���<^�0������L��8��X$zs��x%6&��#	���R�Σ�����v�m�[cd�Ν�^wCB��\�jϡ+)�w������ m�h9p�    IEND�B`�  x�PNG

   IHDR           szz�  ?IDATx��_LSw�y��{����A,JS��� e�d"����z   JK��?�R�X�Q���M![@E�"�a�	�̘Y��mq��'Ͳ�}vu/{���%1�In���M��|Ϲ��_P��h��/.~ō���\����Z�;�����FFF����d��y���n����>��G=z�Ç����2K_/1=5�����277˃�<y����u�{t�tc�Z���O&�������^�&�	~Y~���"W�^!8&�
n������XX���˗93r�#������$(0����g�TTT$�=���ο�E���(�B9��������vu�PVV���I?�^^_7��~����@�bQ)Iܴ�[�f� z;ܴ7;�M8\��8Ek���α�ctj�q8��T�+�\�C��cmh�`]:�gs�Z7Ji6�8چը��F��T��_ M.�u/㔆c�7�T*Ł���#��f�am�S��QSkB�of�	���k���",,�������T���h<D[��!;��nmE��P.�j9]�uz�R��+�f��6z��ilS$���pI��(r6�hs�� ��W@�P�EJ#h*/D���ݹ;)��%9y3�����Onv&~0HLL��g�v�Z��Q��:�nM�-��� ���)���n���d2q�p{z*�q뱘�dlO��H�Q�*rr��x{[*���������;g���vj�����h��t�Hx�Mr�w�;�CBB��e��V��K�[T��t/	�$�!�05=}���0�@�����&|Z�{���C=ty���N���E4U�p����gff�c��8qr����w2)).�ek��gE�y�T%��&� ���mIebr�QaD�?��T��`G�ܸ��	+Z�xi(�veSu`?--6a�!�\��h/u�MM���CZZj�,,���R,�:�lNJ|Z�W>?�a}7t����R^�"%%�(�X��uw�Vs�D��q�j�DDD�-��`4��`%h5-Y�q�W)+)��P)�<��z��u�Z�z����L�ӷ��V�V���*	��WG���Ќ���))I��Mz   ��_Wo��t�oϋ�	�k�1���    IEND�B`�  ��PNG

   IHDR           szz�  [IDATx��[L�gǽ�՜[��0J�P�a���������'h�(J�Ж
=�
EDA����\69��:�v��m2�x��3���˲������0�$K�$�͛������=�����c����?r���\�r���Ŝ���~�����̓{����5n]���:���<{6��'O��}��>�����'� N��S��=ϣ_~ejj�������{4k��Q\�������/.�������S&&&�x�"M�������/^�ƍ/��.��t��p��]�����@����{;�d�K��0<r���{�.�̣G�G�S����JP 4ͫ}�-45�������� ǚ����Ĳ+����:�
�M~����Ÿ|U?�NeuN��6�8{��=A����j2RpȄ���B���	�ϋ����H�6s� ڎV�*�PXx�"����F�KJqy�ԉ���g�#x �k�?��Q�Xp`� `2[���[�D��<�ݙ[)w�p���́�pފ��������9�#,,l�#BgU\"��H��ӊ�h`�捨�
�hĂ�t���(�KMحFBCC��
���`�+{;�Z�mM#{�bc��ܞFl�Zҵ[�x�ų�D�E,_.eɒ7�[�Y�~ZM�P���<N��l޴u�Jxf�ŇǇ	��ݗONNn\���q��U�� �j�����'�8���u�DBBBX�`��E��Dk+UUU/�������USS霱�`rq�8""�Ѧ��](�i�����9Z���H��+��\�/)�իW�����]��R�33�e�/��s��/I�R�%�'�>�^��x �
�}����g��~��Z�g��ŧ^����zFFGk�����z�t;���!�>��T��H�Rl*ǛصsY[$�곱Y��r�gV�.V��B.�a����PƺDyz   ����䂪V��L����$&&�o����iw�oA7�v��| �)A�������1'�[�rd1�PVb���+W ��a۶*��:@����5�d���&���9���8��47$'g�Lƙ�����
Bs�qn D"Q�T�B�@�0�SR�l�ֹ�?f+�]rS��    IEND�B`�  ��PNG

   IHDR           szz�  �IDATx��kL�e�g��&F� C�\PV�w�k�"RXK鸴�0���^��!nܗ�Kt�Õ���q����?�f"Ù̌�O��e�$&�����������yΑ#��}��[�1?����ᧇ*���-�m|���9�ߺ�)�wn߁���A��B�8���#�����Ǐ�p�!6�n`ueCCC�@����@?��V������}<y�l?@υ(��mZff�����k�簲�f;�D|}}7�n�ҥ~�� ����m����azzږ�Ų���-���q� JK˃?��L������119�d�>?�v��> �X���	�=]AՉ��a��]�yʌS�$�3���Տ胸�e@��J����x`��&��j��R)�Ѫ�(/����B�Z]3�j���DTCk+��{CW]I@�G�X���s�8W�@�V�����л:�^UG�H���VR�z46���2y�2��Z��]PYq�>���؈��b�5*�u��kiGK[�I�R)D.�P")����w������WAR����p������_�����FLt8
����K��$˲�<;k~�@�G����]/�3\�x�$�9)HINDlt��c!++��'5��2888T?��y2E�AQ�����LwdDG�/�H�f�B$̇�M�11��⧁u�i/x���eM&�>�����\."Ã��� >.
��j�SR�m�;ZѨ�CPP �����;d�\��P֞EQ�({{{{r�QS%�X��L>��шE + ��r����z   � ����\��el��:��ѿ�<;;;??�<=��9;;��#G�^�� O��<���'-���e�SծM�bٱ�W��_�#�ښ��b��!(=s�g���g�ڄ��!����e4�@&$M���;���&����� ����W�.#�鲇-	���d2�^a�����!:&!���HD��!�����8��-��1��'�����f!�b�{�_�kl�N��������A~>q	U�2���P������J�M�?��20�|Ȃ��=���������*��@�(�t2��b����z���C)?E������,>-Z(j��'����TZz8}����S||�3�(.�����k���Eş׍��]њ�    IEND�B`�  ��PNG

   IHDR           szz�  sIDATx��[L�e�IL$&F	c�:�)��Ph�Pl�a[Z*�+k����
=PE$�&&r�	x1�rư�Ɍ'��#�c2`w�+���+�		�%������=��>����{V�}����O,��X���>�Ə����}l�����O����fs�� ����vvv������-<�|���AP.n����vcss����'� ��,�}wan~++˸����f����x=����6��<V����ֿ]���/XZ^Ƅ�E�[J%�����o�ĸk��������GXX���n���N�Ѡ#W05�	�����p���9�1bc����K��AL�^�ؐ='�&t۝h7� ���@ ���@g��: U��KP(���P6�`�耶U�^g/���0���p����C,�@Z� }�m�&�DD��|�N@G`(���6���+x[�G��24Z��z���&u yyy���T��C��X��sW��_[j�B�h��O��_������!%	N�����A0��PR�F|�ia8C�@)iAMe�,&�U`rj��e��� �Ț�=�5�����,�D6�����8��z   <�fe�s�QXp!!!n{<���É�����Ƣ��"^4��'�(��������ע�d ?��s�հ�<^/�ج�É��ML`���� ���9RRxHLx�FmZ�#�����^��vX������ $�Y��C�Q���<�υ�RX�xp8	HNN��� ��"����	���:�m���1?5q8v
ee��R���{��W��Y\Z�^���a;�u�s��X]���^הR|){�o��)�=믱a5�Vk%yవ�J9�
��a�&��N�N������R�r��<ݐ?�`Z(|��Y�[?!�&#���j���2�ϳʊr���H$�p:�Y�������n�6߲�,�Ĳ�����i ��qq�x�緳23������Y����闡�RL�#*���E�H����k��,&	d&驈�=����D�t:ʅ�>��|�)��c�/P�U۲z)�rsH�7���\���2�E8���+%����J��m&����87��=���Y���ь���    IEND�B`�  ��PNG

   IHDR           szz�  |IDATx��kLSg�1q��6��\�Vnr)іb(�R�b����B/��\�0�؆\�.�L1�X��"k	eͦ�L�c¦�!��a����6͖�pH��INr�s�����y��=��x��T*��vǶ
���������K��|o.�"�|w���m��gX��>��~���c\��:V�`pp���u�bbb��������ڬ��e:ZlZ1?����\���7���	VWV0vi#����055���p8�Xp��n�Z����ڠ@&�1���4����A_.����ƷX%)p8?C�N� D"��@o+�C`��>Rt�_��ǟL���p$_��h&�>�����@kh����ζAo4"33III0[�0���hP�5��P�P�jҢ����:t�ݍn?�PJ� ����QVz   &F�P��@@��GLz=���
�j�>��.Z4JXZ���7�H
���&m3,I�T�#�����Z\|�� x\�Q�@{��YRf��w�j�P'��XH0T�������w�cddx�.	��o��׼_�Jq9�
 3$Y���C(ȃ���Ś}���sW�y�jKڶ�������D`�^7����q���!==�I�8y\;�ρ���_f�p8#�#�67�����M�GFE�@D ���!��Zu8��9��ztwu�@J"�2ӈ+�x.��1;d���۞��vz2���(*�#=5�P+�d�g 1������>u��)���|Adrr�r9l��7���|�)�D���UbDGG�YRBl�GllX�������� ~��h�~YMf��������AFF>��2�2v�� "�����3-����6I	��:J�/e'������D�#�H�'46�ގC&�l��b�G� ����tb�
u#�Z�[��D��s�ĽX�6*`�)!.�F0A7i?���/,�Ce���l���bH��0�oYu�l1��@oo��f�� �e��zy��C&��b2V[#�A��4��JRI�9P�U��Axx�-6&�� woHH�����/h�=����rQ8Q�D�9����ږ���i*�"�� ���Y)���]�\2����J�R�1>nǩ���le��%�Z==�    IEND�B`�  ��PNG

   IHDR           szz�  }IDATx��]L�gǽ�&~ⴔZEǗ~ԉ�@"뇂�Ph�BiK���+��LT�A\�fS�Q�
�ͨ�Pg4x1H2]��r���1�Y��K�d'y.����y���w�rh�k�=iϩ�FGF�s�C���y�[�޹˸���9�o���GÌ�<���<��!�ǎ�����ĉOy��3^���:;;)**R�
p���k׾��ŋ^����7}<ʃ��<J��q��{�_��z   �+�W���k׹!@<��	_�;GgW�x &�)���nz��r��e>no�HG� 2��{�짡�A<����)m����*=Fk[-����=á�CXm6R�F��v� �6�}��Ӊo�v6�a{MQQQ,_��ٌ��%@Uy	�5v<n'v�g�o���wo3͒��v� ���7j��t�4lDyy� ��S�eW�lv�x ->7.��&��RLef�u^��j��R).ҋ�*z���[�.���R^iǷ���J�fr�-��r�?�2080v�T!dA�̘1�!�ؘ(�͝C�ʕ�OK#;+��U�di��d�M�٩��677� %%�0�`̟�\y�R�[2ѨU(�������%fQ�_+@��[���驫���[򤤤���(Be�f3G����2�HO_+H�Ⱦ�����A��JrR<�fͺ��;���c�~j�>"<��ձ��X��@��XˋIP��V��d4�z��D¤I�2_}��Rd{u�ؓ�Q���!�6�Ӊ�\������h���`�p���;�Iy��Q��'H�_O��NS``�T*�^��w�ĉ���H�,%""��B=����I�x�?mo�ܖ͂9��n�DIֺ,(���gNaO��ۥ�����-_��:��O4O�ٴ��5����HOK�H.E�+�xw��"l9���G4 �AOV��b1���Tl3P��e�L��>,��YZj
y�Q���)�䒫�f"\ܯ��6�
;�܂RY���<��%K��Y���LXP&�'HNr�i
����^���Ӑ�eD�.HUؔ�|t���b��Y�Ř�>c���_ZnH��D��4�&O�|`�ԩ'%��C2Y�3�T���>!!�i��llv;wxغ5K���"T�����,:�Ge|���lJJ���x��'���U��    IEND�B`�  ��PNG

   IHDR           szz�  PIDATx��[L�wƽٲ�f�aNDE\WP��Z)�rȠ� �E98i����Rz   )��0a2����]�Wn�FL�'�b&�Z�K~�$Y�d.����ɞ���{~y�������|z`��`Ѕ����R�ύ��>�`�[�����]�\������h4���'��0��,s���Cn�ܘ���Gt��7###ܿ����ѯ����DW^�OT���&'�b��E&/]����<mǽ�14<�����U;ř3c\�r��SW�Ifff������q�	P����v�M\����A�e��u�|7����f�x Z��������x�b�(]==t:ĉ�'�l�0���H��|�x��=�l�d��j�˞�f��l��C&�Q먥��I< ���QO��NEeF�U0l�L��};m��8�e��8�d�?d۶�ss1۪�2���l�[-��,d�n�x ��pX�;j(�W��4R[W��΁�ڎE�I��m��/�a�����V���p��އ�T��PI�����I$q �R)^��R����8V,dY�Rd�l��B��BJ���\|||^,�J�j\���;���A�:��D_�<��J�l�$!%9��ʝ���>��s��3������jA��%�1��J������K��yl��HNT����L�ѓ'������2_�ȇ��l�.!|�b�f=
Eq�X��o��k��ʸ5>r����k���~�������?�Ѥ��NCKcM�1Y�:���=��	}���//���D��A�{������^FDD������a�bɍ�bJ�b�d��E�tְ��� �GG1[,�L����=vd�`!��LO��O7�M~�S��g[��(,����g9䒝�I�� ��Tz;[ikoaM@@�t��u�UQo�ZMYY)1�,-nB��%�1ˉ�x}�x��TT������l�,G��B'�$%ŋ>�)�����XlL=����X,�KD7/))yӐ�<n����B��7ii��8��w��t����V��5k��d���Oȿ�RAfF:�k�wBAjJ��*D��<�B����f\�Z���9Hz9z   ��K^��6��ER*̂�l$4�����WQ�|����    IEND�B`�  x�PNG

   IHDR           szz�  ?IDATx��YL�W�Mn�6�҈LӲ*�"�32T�Ev��Yؑm�EY�B�qK;\8�`Հ�bS�Zқ�6�����]����Uo�Ą�Ĥ_�_�7�{����oÆ��SS?�9����º6^Z�����|r�S|� �%w>�CO��j] ��������Ͽ���2�\�pɛ��u�r]���/x���3�<y��������?H
`wL2e��`aq�������/>甓�wG�Ua~~��ׯr��5ffg����awpkiI -p��9� *++�ό�dN@\���5�b����6_޻'Ը���[: ����Po����x�����0>1���,��m[Yh��h�ޱ^��:hlm�o�8mt�lh�ZzlV:�:�(?���@ufM�T�hhl����.k���ʐ�ԑ6��s��˧B_MIi� i����#~��$�b1J0:dc�����faA�:=Uz���T��Ds���"���P*���@�`�5`�9ʠ8���~�ZZ�5Q)�֕����
�V��^777����N'*2��7�귅�����'h�V��:�[̈́���-�\.����U�5��Ø��"U�D�|U�b2cd��D29~��S����~�� >�^����XCj�^��R0�VSkб;)��!��(Е�y���}BB��]�����bB�P��L�׉F�A\l	�h<<<شiSٚ{���-v�6��(��Zv�#?� �]m���C�J���}�֘������x3����ظq��u ��zoD ��U�d�#��y��������Vi))���G&����Ixx8�&�vb�*f�\��kS�N8��?���g/3:6��b!C������Ҵ&��IN��Ŕ�ƙ�J��iȓM��b�n�l2a������$��gO�H�d��ߤ��*F2;�l�1�3-��|�<:Ez   �!-��!��^I�~6+w�Xj�(/�CIv���u�kU�פ�QΡ�l|�mx+*R��}�Q2q�qZZ�Z��[��R�Qё45ZD:*I���$RQR�ܼ����Ԋ4܍\Kbb<�Ѱn6xzz�Tg6P��E��&::��׋V�=s{&��     IEND�B`�  c�PNG

   IHDR           szz�  *IDATx��[L�u�I�mo:�23���2�6`PHǸL�ri�r-��B��P
��0�ld�Lf"0l���P���t��h����_�|�?�O�>��9�s�����*���j��w���c��]��ǣ�-�����=Xgdd�������cuy���=�N����_���Svv~�ɯ����-���c��"���LO�`~�+?~��/y��9;�;LLLP[���k�ɗ��feu��lm��������0��� 1ϥ˗�15���`c� ����x *�ꍉ�!���������M�~��_���c�W��;�|����h�v3�F�;������o`���ݔć�On������܄Vo���Aw� �mm��:�w��\UI��U<��B�ˋ���Q�������@�V���F[L�� ���qZ�����Ց�����@}C��0V���iqwwG.�7�9�P���;-�Ft�&J�5��+)�h���Q�((/U����� _<<<��j�⹵�D]�I�B� �.�B+rs�H��Q! ��2��8-�0����m�Ef2��g��#��D��h_N���amdb��{zz�b:+'""��"%����`N�e��&$( SC5c}x{{�=��07�p22��jc�HO;KTT��A����.��J��L���1,&���dff���"((� ? �<E^^^�$|��'ve�c>����q�e1H$o�{�����Tt8�2�:ACC=9�l2#�x�]���D"1"$?'��#��^,\"+#�����}������>G����#���z   �_�񵙙١�[��r�
#cc©�HOO.�������ͳ�j%z��V������'�t:��Ԑ��FFj2��L��<*ԅ8ڬ�{R��/�ZM��T���\x����Q�*Of6�_�ƴO:��N���,����8�(((8�o�K	&>ԗ���ݽ),���X�U%����D�'&��.܂�]&%%bk�`28t��� �-Fd�DG�P��si��+����/-8x𠟷�׏'#����H���0:"X4Kn�ǫشnmgLp]    IEND�B`�     #�PNG

   IHDR           szz�  �IDATx���OSw�K拽���2J�3j���6Q��l��A`@[�R�-e��>A˥�Њ�]�2*.��e�D�Ӹi�3��$C���&�/�5Y�Innnnr>��9'�ޔ��k���񇇃~�I
�(��r}��K����{�{��~�a	g'&���իW���#��e����ˋ����}��σv8I����...bmm+V���GX�_�?@E��K� Q_��s��D"�~�L�&p��%,/��3�Qh�z����0��8fgg��3�{�6�Z���7�ř�i�z=�
:􈝍an�k��.��B�u��.\���|>���Z�8HD�Q��Lcj�s|v.�O"��i낡�@� ��ԨT��mp9{0tď���X�lP�����x>�r9:����h����~�I��t-�	�~4���R
� ���t����uu��X��	||beee�-z
�}$��6x6hZ�(�Dm-I<||p5!55U�ת!�J0���a��JeM����R)��"���=}lv�d0~�iU)����IJa5R�!r%%��� ��|B �tde����豴�����{s�	�P*���ڲ��
�:qb$�������I��@�fۛ��0c߾=0���h�_�݈б u��D�rؿ%n
�鑓���y��I�/�vvb4�4j���f��Ҏ�Nz   ��	E��De�4$_�;�oo76lxL&��v@V�E�yЊ
p�ͭTި**��j5�bb�Tr%�E�^�}=iB���,�F^	�A���,0��,���^�g��d")Uہ��
�a��QSߐH.w22X?�H��T��6x{�`��ڌ��a���������w��b��Drg�>�"'� 4��eE\J��
�&&}'�\D\���؉��t�5��[�?T@}�j��1-xm'�x���+밽{vS+�BA	�b�b�y���2�oP���v��~�B�=��4�F�_;L4\�A�8    IEND�B`�  �PNG

   IHDR           szz�  �IDATx���O[uǹq�2��6Z��		�0�Ȑ��xshYKKyiK���ʀ-0�Dc��gHƜ��h�4ۍ6�H6��K�`LF�M�_�Cb�'�]�s����}����_@��9�=�8�ͶkGE���^�cu���u����{+wY��&����;p���?���K��ܸ~���Gܻ�3;055ɝ�����M���c���q�=TT�R�*��T3�ٌo�ZZ���4׿���Շx��4��uA[��	]���̌����J��/��ƅO/��`672'����.WgG��}k�o�]c|bW�� �n� _\�"80���%��g������,.@vV&55�8v��vF�����382����h4�����)**D�T�b���n��i�l7��*��0��|2�>j��*U	j���c��h1�Q�,��T�E���IMM���nF�P�c5	�4N+jM5�F3��?����{��{o ɋ�5��j)*:��H?î3�t�+��`���lF�ѡF���J%(JN�d�R��ű�����P�����Y�/N	��^���F� Ig^&�3�aR�f��R�u��j�Vk�`K̠�!��@��	�P_EKS�н45j��j%9� :aR�:[��B�i�ҷ�#6&�w�h6��|	�݂��D||����l�z   �@��B��E"	!1*��=��A���BJ�����gDp��J�cN��ݻ��%��(���i�O�T�F^R�%%*��&ϟ�?��\��,�۷�=.�Z��2t�|HBB���6�	�w���þ�AAAG�JN��ӭ洘��(��'>!�LR�P�@~$ݗ44T��?��S��eN�N8��da���7�3d2�/�\�An^_N��z���SS�I���/�%/�Hġ9.t����	�I�"??w]�K��D֒C����Ű]"�#;K.�	�&�@��a8�����V[��P��i�xO����(\}��    IEND�B`�  ��PNG

   IHDR           szz�  �IDATx��[L�e�wg�0���s kȄ0`���F`0dci;�ʙBO�P�J�ˡ[�F��`#�`/��h`�Ƣ�7,��.��a���k/�K̞�/�y��<��}��ݱ�i��xp�ã�M��Zd��;|���LOO��q��x�Y囥[�Z\���G����- ���XYY��������~��s��Z�������L^�dff�����߼����Y�Yx>��j�
ť�LMM1'����>��c}�W���p]������Y�n7�A'�������w��q�p���+.@~��A� sssLL\e~�>�t���I��.L�-�?��^��l1�c?ψˉ��������lm���SVZ�N���˂�d�i�D��Ҩ�P[[-���	d29U%s��ʛ�����5(+�0���Go/����DAa�V-f�{����r�Q[0��#;+�Vm-2����NF�}X�Z�+j��S�P(���w�h&��{��&3�5��*2�_%;#��G#?}����(,P�S������{CC���b-ȥ��@��p�mFڅvt�3SS[Eey�_[`m�%+3�]KЩ�i1��	����S����#��Iڬ歯� ���ԡ!�B�C���ni��Y��t?���%��z�FUE{���z   ��H$��j����y+mFE<��!;w�C��2$::��A;���	��S�J���N%IIM=Va��Y�pZ#��~�x�r�o%hk�
~07�	��{?pс�I�6$%������K4�j��^��NI����3�> ?�]�e�3�[�p(֗4ⅰ;�/�0>��������;(���k_���=�� ���>��<ee%,~1O�`@�0b��z�99o8���Ě�;��ʼlzu�d'Jqgee�>K̿<"j(_���"�ꌸǂ�~~����H9v�s]��9�����L(��O��Oχ���S�����Z    IEND�B`�  ��PNG

   IHDR           szz�  �IDATx��YL\Uƛ�#-�(jYf��2�Դ�����h� S:�t��m��e6�2-�@i(���b[�Q�_�1Q��֐4R�������>�LL���{Or�������=۶=ѿ�7�K<��w�o/���
_�3sk�-1w��x�v�'�����W�<z��_�o@Ss+++,�>~���:���`���𩹹�<�?���ɫ,.,2+�>{�S��e�����m
��J������fdh��;wx��W����^z��|�V��v�W�\���55~�������봶�� ==wG;�OM16>ʍ177˻��t��`w�|`�a�Z�p��u��ɱ~��/RS_������jQ+唔���Q�/�R��ш�hF������())�t*rrrhsY1���@��G�T��}�nm ��a�d���դ�b��nn�XZ:
e.��g}p��9RS(��
 Y�����X&$P�F�%33��7��Y]�����I�%9�G�x��~�Ri?_��0�7	���ij����H$�X��:̜�ECm%��r�-��s�h��x�f)_���& ��h'��|*ME4G�Ҩ��a">>���7)+-�>�ɠ�)*><,�����H;B���tg=	�DD��T�L��}���<EAz   ����	

$R��Z�a�wل���"-M�?��� 2�������蹖��Q��:� ��d����8����/>�`<�u���曍�w�Q�ɒe�ȑa�(C"ߘ�qX���x?�2{�"�hGIa�#��K4h���=-#$d�F���%,�� *��3�šs�?=9H�AGq�
�:����O<���<߃g�^�H� Ǐ��P�����i�V�gg` �^����ߵb���ў}�����n��z)�(��[�S�M��S�ș������-yK bcc�����J��🪪2���D�8�� x���|����'k!-n    IEND�B`�  $�PNG

   IHDR           szz�  �IDATx���OSw�y1Bdji��/@E&,vD�ril���
J[�Bo�����B�tm���\Dġf��tKt��\��m�M�#
l3�]�gg]�_��d��7''��<����Γ_X��y�dU�999��\���w���~_[ǯ˿`i�1q����<z�����c��OX���7B`n#p�{�zn����'X^Y��@?|�|�BL��`?�\ŭ�����ݾ���?`r�:z?�@�T��#���/�уX}���g�"߇/]���Z�k��p󓛘�N����"��S���x���8���N'&�q��4n�\��Ca�Z����IO��7���q��t��h?.��aiCO��Z���q�2Y#��F��z�q;�"φZ��D"�`zr��oܑ7ԠV\�!��V=��r���� ��oG||<_�,CYy9<.3\#�D+��2��������:���т|+*p�˂��n��J�՟@C��5�'��{�~����`�Y0�(���A.�ge@$��eo�T*�@ �:�����}�O#v�V�wl���V��%�h��`3���i�����)�1����'������\z-����UK`k��P�[��y��4�0(N,���`��`�X�z   G��4��هvR�J��{wJ Q�0� M�RϹ�.DFF�.� {Wڌjx�L�;��R٨}O�O?%��*@������jtbccǒ��9��M��D���JNN`��sCR[�tN���v:������\��C�X�6;���r ��~�[ࣤ�G��T�4K #��^,����mq�c~�� ��㿚��{��ΝI�hr8��tr4���ҰeK4۲������� @ffl63"""02�V%A4-
�p����*f2�?���;�#>��r6�ۑ�DGQ��/�;Ȝ;�:�d26�v�$����[1�W�&���s7i4ZJj�ِ p��6ZZTHJJ�&�弜 �?��ݓ�mK    IEND�B`�  ^�PNG

   IHDR           szz�  %IDATx���OSg�I���d2`��Lx���	�¢Ek*FM]�JYK)���RZ(�J[�RT���B�/qq�%,1S���,f�Ncq�N�eٲ,~���zI�x~�7�7��s��y�=7"���@�1�������].W������[<��>V>�zp��=�ڃUl�xG��O����V�ĝ[���(����:�^G9�Fۈ�׮b�������[F0������!j]0�n�1,|�������sp8�������8���Z ��t�;2���QLLL��`}-���e̜	`��CEE�[�TUU��������	������o�v�K\�����L�J ��o7���۱0?���K�%��@ ��1�	���B�J�ʩW�P]-����لKgN�7��jE��	.�E�8������|�X+���.��ܽ����焢V�N����XJ f������i��Br�(���1��E�A�����a4�Rw
�'�B�����#G0����`V3qDu��lK5 ���m>�������@,�U�����R��Ґ�P�˩跙�ϝ�yy����A��خ�CP̃��]�#b���w�0����GYY����hP�Kz   X�.� �&%l��pv�b߾�h1���BGK��LA("22�J��-Mu�<��f��mM(��O rѬk?�Q�&Ƽ(**�X��;s����=��7�ì++��ի�W��/^
+@#�`vr�����x|3�6=�_K���R܌d�3�P-�E�ax7i[�	�9l�H�o�S �섌����x�MGƮ��л�	�\�߆��l���L@N��\ ��"r
T2d�г-�/���AIIqx�����bbb�II�0��l�Ԓh�^[���d�h�+7��p����RSS�h�W�c��aR�:�,zt[[H����#(k�6Ksh��333�QJ��q7�er_�T ��2���8z���L�`�A�K�nd�`0�l:��^�@ȧ~2NHH �q0�;��m�NÁ����z�r �H���|��OҘ�T���/HLLܓ����s��Y�!�g#7�K���    IEND�B`�  8�PNG

   IHDR           szz�  �IDATx���O�U�IH�^�:�P��&-��Q�}	�����B[��(B)-�e+�*��b�l�m0l�u�ƘK.�M�����l�l2L�K���ך�/��d�չ:��<�{���������������]\�4��U�������=���&6��`gc�b�p:�@j�����1�x�ۛ[�gk֞�U��gTXZZ£��r���{�D"����w�Km
��!��]�չY���O���z��!L\��B�Ȥ�h6��.�afv�SS�n�>��6��������@�F�R�	�qg�n/܂�n�Fd�WV���@^�*U��2 �X\��Ԣ` ���ؿ���7���0Y,���bQZ���P6)10���z�CӸ��0���p�� ����ܼE&���I�
����~���9���a�h4���FCC�)J >�@�V���r9<�p�灱�j�(����d��z��+S��`0@.��PT��;|�>��Ԉ	�k;�pک�cg��z   _\�BV�
ǋ� ��ԩ��゘��%"�J�mSQ0�q/n^��q�OM�բ�����υ��
V����B(�"����|�d2���*Ι���v6���8�nD��^=�c�i5�p8̘��>1$&&z%� ���K�-�!)e�Z����t-X��H$�mN� �[�✀ݪ��\'
�9���$�ˆOZ��+��pNd6x� iJF���|+��6��\�B�z���� ���}�d�IGv��P���$��L�8'�ܻ���2���!��ǹ�� �k	!���fE=��Y���^�G ;����ĸ7�g�������M���Kw;����#V�|>��i��9Y���.8z�����(�oP��X���x((ȇRF m�>x����FKGi))))Ԧ@���e��)-��S3;t(o��O��{�z��ɘ�:A�.���̎���Z1��X)��*���M��g ��B�z�w�_Urr23Ṟ+N�;Me��T    IEND�B`�  7�PNG

   IHDR           szz�  �IDATx���O[u�I|��i����V���PG����-̖�t@��)+����(,��vq��E�e��7.��[4&*l�}����Lόɞ�8''���\~�yNT��ռ^�܏����k7055��Pſ��9�����&v���ޯ�xpE��m�Ķ�Alܽ���>����պE9�V��µ|�՝��]��f��p��R���������*._���w����0~�؂���9���G@���<��|><��u�3������:�Wᙘ�V��P@�k������"�V?���N ��E�riy	�cgQYYi����P�˅@ �Y�e�� �"�f2A"��Q�z4Z-��X:p�������[�
���a.��Gzz�Ͷ�j����{��Qg/�P����h�J������/�*�P�Up:,��q�ـ�z   j
� M
>��t��I��W|���Q���X��^+F�l06 ��P����J���cyiJ��Q$����#����dD��e�QW������B�R����`65�d4���\�J�a�h�`��|r
���8��K�f�D"��t�j�Ao,��l��b8^9�.K��d�*d���ay�C��s�kY��"nj������<���RS��p����u�^q�9�ɀA�E7)��L���&dfƳ4�휜ltiJ#��bࣕk�UhÎ��E�B-GOF*���������w$'+�#��BR5��,���P���yJs��� ?��"��-���O<����"_Ϲa��!>���of�#
�)W�E�L�WyN�P)����ֱ�9L_����n(219r��Po��=ԃ��s�]F$v��w	II��p� ��:�a
̈́9�ydy111�Bd�xx9-)\V�3h������J�{���`��Ȍg�d^�LzX��`�^���G�P	���Q�(,�%Ҍ?;�a!�`,J�e���B��������XJJ2�����c��_�FK>t(�ӨG�����	�H7n�G�    IEND�B`�  F�PNG

   IHDR           szz�  IDATx��kLSg���dl]�Ep��ґ�Ea:�8W)J�����vPZʠXn�pF�-+((2Z�CAT6f�l�̩cW�es3�c΅-�_��o����,�9��I��������_��v����C���w�Xk*~���X������D�/�~���&��W@��qg~�o�¯K���?a�����Ƞǥ�i|�;�E@��y���p{�8��C��F�3�v�~�9��	8,,,������TN EQ=��]�!o?����=|���9�9�~����6 �^�98t�I?������'׮ctl����XK�D"I����no���8�>���y���t_OQ���~�6����'̦��磵�6[-�Nyq��(z   ���sB�RqiOMM]"�����.���L��c?��t��儩��ټ���}P��(Ԫ�P)�lyG;a�4���~f��|~�o��95rz J���Jsr��dE_��uUP(U(-+GsK=>0D��M�A$!�� �L�j���u����j����EyY= w.3�P([M�J
!�J�Z���r-6df�!��H}%.
�p:���M�4��b�ݐO �`�㠐K�n�.|6{S��b��59	�2=�ײ`)-D�Ռ���`�<�MI��(kR@:k1sy?��^��ɨ�u�J����ּ�����Fp��``����)��rz��QJ\$Y<Xօ�}�u�L�w$ 88�e��^Z`
�*�{ׯ��d2�'�=�9���C���T6\mT�ʷy�͎�98��6n|��*��_���)�&S�앣���l�z��)����q�L��Qd2Ӡ�����AsC5Db� 1l����Ih4�����{'�9|��ހ��lI�?R�5`2���(1jp�`+bc��X�DL���BDDDT�3x`E>�͛7�X�c&&r��&�M/����oh��L*Yu�����n�����]�(�H&WT�6�<4������$,�ǽ��%)d�z\��_��hA���    IEND�B`�  7�PNG

   IHDR           szz�  �IDATx��}L�u�ٴ��Lf�P���P�dPg� �;��!����;<���T��a��œ�P���dv��4P���yP2��@�t2e�bkM�W?����s��������������4k�u��*�����=3̃��ܟ�cn�.wo�2w��ż��������͙ܘ�a�Ͽx��?h4�u������pu�'>z���4���tww���,n
V�ի�����^�31~��3��L�����6qvZ�:t�t:�:�ɵ�If�������9�������E��L����#���wRXX��?n0��4'O�����^$@R��^Yz   UAKKN``�����q��c�������=��Wa4�������oz���`+��=���%99Y����@��읓�B�Z�}�����>��Ƞ��ĂN�#55�%Q N~� �V�EVv�M�Ԗ[(���Qh@.W`��-t�����###�>yRM�v�lB
Vὅ�\5�R}ߑN��B&��I�.i���ה��Q�Q�%/O�V�A�S����?������X,�����m)D����J�2AH�D��HLLt-�*7�Ag�~��|�Dxx8�)I�w��Ϥ�f�|��}�ڐ���r�ܵ �z��
&����������Ǚ��0`�U�\�֯����:����w�lm`��E�_���p�����HJ�oc�/�e$$$��˟C"���M��Z��s��>3%����ޞ�~A���b��BّA��^˞%W�Z�O�����۷~�`0���%H��#E�M�F��q�u,���_8��NP�b�<,��?�/l;^��B��`d	1h�q�-#>>N�U\��W&�P*��Z�2Q�E ��@�0T9*q6�����w'����DGJIM����@wG���߄�viii�Z����h
u�t�9x�ח��z֬��!����k9��o�+P]�^�K7Pl��6P| �BN@@ ��������+V�aO����?���?Z��UAI��m۶> 7�i}=]O��=��$ZC�*��    IEND�B`�  '�PNG

   IHDR           szz�  �IDATx��mL�e��Jlk�l."!Lf��W%4�����v���p� 8<�5� ��;"A�J�i˰���D�U��>d�X�����Է�Ck��t������뾯�7lx�"�n�������֍�X'g�}�6�"^U]u1������?O���̣?�\ SE9w�Ǚ�β�����<V���籜�����ح�����.��q�����!��tS[[+-��V?lniO;@�19����p�>��m���� z   <!@�*���^::;�tq ���1'�a��,5� �`䔥�§���}����##W�?�O�SM&i��mڼt:�u������FSS#�fʌh4���4%j��*���h���\^��Ԉ �|��Mhhؽ���IJJ�\�E�u��%Z�3����r�����E�T�^���1��)����xS� 66���Ji ��:�7?DTT��LRRRh�>��:�2����C�J%F����vvv���F�s���acc�6O���/�## 2<��PLQBz�ں��ϊ�vv���Q���HOTP^�.�
/��A��'����2ry��|T]ɗOo\����`0�j���G0��S��
D������ݻ}(-+Y;c��ζF�����u�ł��DF����*^V��w�d2[�����v �!-��ȸ~�*�S���M�lV���D�|E�𝫢�����խi�E��|3�uv���d���$�^ϑyp��^!�ϝ��'%+B��X�D��a�B����|9�?Ur���BtxY2 {{{A'V��׾C�/�m�+��3<t�,!�UjA�> ����s$&&�y���� ��Ju��':�u�G2}Aqqq��<O��`��z:���� G�!lmm��d��N/���W��B��ɀ����.��O/O�ow[��xc| 5Ḻ���e2���X��z�wC�*Y��dee��h��iY���cf<vy�� 8;oQzyyN<�3�/�/Y�A�W9�    IEND�B`�  1�PNG

   IHDR           szz�  �IDATx��L�e�]3G�6�����	C�C]�䇿NA9���8��N~�%t�"0�����&�4+�Y��f��e  C�ի/l�G����|o��g�����y>���.Y�4�"c�F�i��7>���k���zzz�n�Z����LM3:��_�uf��IE����)>66���$�����Q?F��[Q��!�d�I��]��� {z   {�����'����JMM��U�h�4�n�����sm<b�'��Op�f�dm���t:�:�5�8�POgG3ӓ��M`���Z]-�@LL�O����M�|���P��\��25�u�
�����3�����f;��n��~�J뻘J�0��
�t��:u:����`o�b1SRj^�^_�2��^�B��B�!�4����C(SR���RVV.��D"i��>�T*�Ԩ�!S�J��BI�[$�OF.O�bI����������L-�8u��uU:#S��J�B�n���p777{���.]`�<==HW+�ˢP$ʉ��N��(,�F���4�ip�@nV���z�^��L�����H�d���GYq>Ņ9�� N\�̱�P]Y�+��}���E�3㑃T�P�QPr4�XY4�l$�����9��m��z��#?����Z?�e{0Pd:Bq����0V<�$H�E�Lv\B��4J��5�w�������K���aa?�S^���@�@V�Z�b�2'�ׯw�2Tx��j�%�ݽCyy9.˗!�B�o�6����8�ݿ}��=[^t|+jғ�no��!���y�כ��g��7�nᘹ����G����B���@8�Y'�'"�5d�v/�BC� � �w ��Xn� 55WWWvl�ʮa��ho�'"b��W���Ө�j||�I���H�F��J��|��3�/�������\�N�Ϛ��U�H�ߎg��M�K��m��������C$(wn$(((St�� ����y�3��^^�1:��F�B��8W�&6.�sg���_qvv~��?��2>v?w ��    IEND�B`�  �PNG

   IHDR           szz�  �IDATx��[P�u�}�t̘&�%h��BdY���v�_�V� Qa�&+B "�� BC0�(LQ
F�D��Ĕc��A�Ox�ǆ?M3~g~O������;�wv�z����W�ni��������Ņ�������g��ڏ?��7����g��?fue�x�z   �w�/����:nl���Lo_/�����\��y��S��ja��1η�2���t_��q�C�@?��]�aei��?�y�`����on -=���A������ʍ�a~}�Ɗ�(�^�^� 2BEKK3#�#t\l���,SӷB�p���E����PT�Onn.��B�u��{�:�s]e9�����d2�:���h2�S��(&/;����WTRPTLr������#..���8�秓����d�j���@�N'�D"�`��e�r9�Y(
�ӓ�W�xWWLTT4JU�U�� \�ng��1rrr�O�Mg����J2����_�Z����C+
@{[#sw?B����ZM,�PTa�x{y���Ac}�AGQ*��m�����$Q����8�Ӗ/SU~�I�*���
',L��i���_��n����uB$'�Ө�6�D����d2W�z�	ex(�����!!!��۾j+!/+��@Y�;������a�56&��W(K�o�
��T���h��-�P*�?`����j!�2;��ٍ�����7
uf&ܚ猾n��}��coNI��<�a���d�%�o�I_�u;��8�
��ć��ajj�\���=���K���>EP���ͳ�N�����|63���3�ˎ|TX~x���$��`q?����ܽ�	66�[���"$Ї��0z���􆃸 ���/656�VV��D)H�SQUV���A�����BH�R��͐ٙc���-��9pM����@<�\ō�Є���n�I]�Hl��YX�s��A�||H�jğ�CC�HMKa����n6���IQ��a;3��S��r223��O���_�}2/��    IEND�B`�  !�PNG

   IHDR           szz�  �IDATx��{LSw��� a�c[��2�S�Bx�A�
$�7�@H�PJ���8^����\	"�L���fD![��=��s:!ĸ�l#~v�?�����&��{s�;�|Ϲ��䴩��Õ5��'_][���o���z   Ѐ��'O�w�W��q�[���?���_x& �#Cܿ�+kklh}}���%z��())�5�BY���$�_����"��.~~����Tg�y���O�������P�x�`���!zz{����2si���	�[��~��wn����>7��b@Q ��ߊ�fcTp`n�
����tv�R` >^����:s�݁�'���A:N��t�(&�� !!!�ii)��D��bi2PW[MO{�5�U:�������,���\dy2ڛ�k4�~�GQ|�RUFc�8 ���ۓg��H$4����RoR�������,��ԛ�� L�����	��"##��#���h�T��D�F]^!�e��Þv._�!%E�Y&:M1�IcHIN$��(�Ғ�v�T�������o�����Z�f�V7̹�4��8�F��Jᾚ�}	)����6��͢�hpuu�F���FM�O:ǚj		�KXX� P�x���c\�2�J��8|[ܻ��u��x{�Ҡ�Ip#""��۷QY�r<@WW+�׾����~���]0T���}K��@A�[���NQAVk�c!�+���J��ݻw��Ņ��sb1dE��^_!qqq%��70��8@������Y


ع3��$)�B��œ��_�#��1�����ҌQ��4L�A.���켘�Gv���(ehʔ4����eEz�$J/8��N^^������Q��?�I_��s��wvX�IMM��ח�н�r�i0Wa�m�ySRK���xRi��AAAc��������=�D�{}v}��D��Y})�J�!.>;��׫7���R���qZ�~�N�����QQB�������QI�t�J�6���п=7=�]'c    IEND�B`�  =�PNG

   IHDR           szz�  IDATx��kL�U���Ip��L��F�6¤0&C�t�۸l`��[�S
(�
�n��M`��ӌdޢN��7�5��62cd�4�į��z   �=_�9y���{n�..�W����Z;���pKK˱�_~e��=n,]�֏?s�o���]x( �!������e���W>��o+�YXXDp�&�����X}��յ?Y�~q��Jzzz�� JU��L2:6�����c|��'ܾ}�q�8E�"a���j��^z��3S����ܻ����������!,���������io7s��^�������C`�<�
���ٹYff����/^`dl���ft�:a�"�V�`46a2���dvbKw/����쁀�����X�r9�5z�mz�fNww���'K����T8���2
�Y�T*F��n7R���PJ*rE55�� �J���>"""�3��Pdf�i��l������£T�k(�/�@������\]]_=VQD��4z,����U)�V�9Z\Ln^Β  V���Y"�F��tt�$'�u`�	Q�*4Lۆ������O273����zy�p0c}%o/�u�"��q$��lG��·hom`�v�-b1O��S�U���b���G_H[K-�/�A��a��t�5گ�q6m9��&�:�n���x�cC%!�eH�~��*��j�gdx�M��߹c��[LCm9�g���1k������R�|�{��:��'���ƶg<���@Li�^��̴��bqc�"��'C��ݙ��������s�� OO&�P���P_[���N{�z�J<�T�;=���w8ݼy��+/�b�h��\CEi>u����]�����L�+��e97� XE�H�`�	G�����`���-:�� �@dT�]���i����^�*��w��p��T*u8���<�I{�I<g__���8��Ot������#J&A"����/�"&&�({fHJJ@�հ}��?bAA2�			������АEj����[.����D]4vd�    IEND�B`�     i�PNG

   IHDR           szz�  0IDATx���OSw�]���e�)�=%sU�bz   �cn�B��
(�
�Rhka-E��A:��!J�Aݦ�b7�`��x��<���۲%N�eK��b1!�]�����$7�����9�s~��.X��W��\������d<R��S|����o�����L���w�G"n�X��ܹ������q���LO���=N�>%>D����11>N�� s1;;��w�\�t��������n��E� <=�gbb�ѱQ�\�{�KW�y�U*�\0g�������`y�:��|��\�̙Nܭn� �����?�������92'z����g��X�� ��h���m��v��̜�x�hh���I5*K��;TY����b��R�E���٥�Rdв�\���P<���j�Y,TT�c4�ەOrrY�4rwf����Th����!T�)F�މ<)�|��b!��O+��.C��/�F�E%4�m�y���w��d*�j1��րM8ӷ+�������S�֭[��W�#3��<5��N�5�~}���0&&�B��� J�r���5�ٱm��}��c8!!���^ff����MM�HMM��h��gE�������s��W��&	�o0ym��	�<��з��e�|��r��LFll,cC^��fn2�c@ �.|��^����h(�=x	���d �_0^����d����k�1h!�:O��"���Y�
ݝ'q5;I_�` ����_V��VC���R���j3�N;�u6Z\u�?����ZZ�[�G�8y�����º��uN'-n7.��)�~����Q�A�Sq>U���<�m��im��&�i��H$��2c3��(��d����xv-�uv�-���H��ҥK]>�%91���M�UJ�uX�����x��r�?���l�G�|#�$�������	}":��^u������elx=
9�/,����IE�Z��pX�jrX�j%�-�H_]�&�UVo�� I�OY��X�B�bs�³F�<����YO�
PRl�������'Q�!�xgM(۶�=���р:GEJJ2z   �aDEG�v�j�,Y���x\�?���=Vַ    IEND�B`�  S�PNG

   IHDR           szz�  IDATx��[O\U���*��@/�F��V��P�yJ3`�)�(0�Q�Z�ap�J)Z�A�:��"`L9Ӣxa*֘��h���q���&1�KvVV���������=����6<2���_��ƫ+L��������m֖�Y��kv���h|����x���<����������+�ץ���T3;;���3�s�[++���PXX��d���^bfv���UVWY\\dN�8�~<HBB�t*����9�����.�?���mgbb���/����r�t �Z-=�=��kB�%�g����2SS��wدJ���&��ֶV��j)5���}���bk�a��a��J`���Pd��ˋ�bb$�����ϣ�(���|*K�TZ�(�./7Q�ב��MT���D4)*2S��3�(-/C�L=��i(""ĚJ�.�z���������H'%5sy1�2Fc�h�'��s���
��'�6$�9CR�Zx=���8��šѤqN�Õ���¤MB_1�(,Uf����R���܉?���@��Z�vP�P0?7���2�kKL�����hN*B)�L�y �LF@@ �����*�Wo������un}9���,��A>�)W�͎t��c�l��AZ�<hw��ب��[�"�p8�"((�N��
xx�BS�[C������'��_�K�M�̇O���ۛ�>�;������&����rE4֔q��� i��8����K����z>�B��_��w[�O�����OZr<g==(�Vp�ɽT<�D�6������b��Ն�޼���7�s�a��r\\\dgb�P�����%7;�2�Ǆjk�s���f�YZ8p@)����ϿIrR<1��*�Ŵ�jv�P!~��he��2�b�(����t W;�(ޭ�����
#��΄�F��^r�?H]e�t ���=|�2�|Jz   �����N���Q����;#���z6''c8<,�[(�q��s�����; eFq�HNN�A.���~Ǐ�R�^����؝ܷ����w�?'eDFFp���Q������J����"    IEND�B`�  |�PNG

   IHDR           szz�  CIDATx���O�WƽqN�Ӑ%�!,�2�,:6����@�A��VE�����ʛ��Ρ$�J�7���s�	-�7�Y�	&�l����>�����ɾ��s�|�7�<�Y��e��/����v�}Ê
�2��$?����'K8�p�/�"�ǎ������s�=}�?��{�~��G��Qk�1==�s����,׿�p���@�V�M����dt�����]���dvn���K_%#3S�.���?���da~�3=�]��L7n��޽.�؋����%���˵���i&�&�`n߾�ŋ}\8V<���#���=�9---X*-���311N{{�[[8�T-����VKHHee%��u���PW]N��(���5�1�MX,&t����R�����|�Z< � �c3%:�hT��ƒ�����jlf=Vc1�����T���Pc.�l�`4Vp�H>�R-�UT�����U4������V���ŁHS(8|�]>��V$��N�\.g_b���s/��y���l���e2QQQ,�111DGG�����:3����M�R)2�^�9�8u��˃}��\all��%Zf�N1���S7�s.xCpp 悼�<Po����Ip�F��~m-w�L26r�o����P?�C�ر�z�'B,շz��׏��*�;�9}����7q���q�����9I��S������?���~�Q �EK�k�1Z�h�9�a���p�N��v����֭[際[�Q�ǿ<��r/��@���5�cwc[���V;͍V:��45T���v��h��{}��	���9��EI��J��T�Jh��P_]F@@��_���縐z   x�k///UF�E�~��U�]-���*����r���=`0+�8w����R�����Ir	�2)E��b��b7�����(���������ԓ�m�{$ɥ$,C��
�'
0�Tf�k����偁�
����;�g��d1h5ˊ�Ś�2��tE�C&���q�&�lق�ߛ|�Czz�� ����R*�P�
�OD�.���̠[ i����}���HJ����B��]B'�ԫ�����U*���B    IEND�B`�  g�PNG

   IHDR           szz�  .IDATx���O�gǽq�M�%�.�Pu1�3-�sʩV��&:F)��`)H[�-��Y��0���8i� �z�l�8�m�n�-���������yo������Â�s��<v������Ǘϫ�o�>���яy��C�&��;>ż�[��͏?��Ͽ0�t������{���\�xAz��N'^����In3�����M��ۋ�j�L�Y_���+=^/��S���0>1��ۜ;w���ϑ��$�&����A&&&9����S�������Ù3=��{� �))B�4>����[0$�:::�}��.:?�T:��)(9���Emm-%%%t������p����ZZ��������r!n���cA>fsU����jv	DXm6�
�y���h��d��O��!���L� ���(z5��Bnv[�J�2R1�I琣�p���/@f��>�v36�M�����Ņ���Q��$��d ��RSu$$$���H5���˾��ht-m'��d��j���ܿw�H�;+e�ީ��~����z�E&�	�J�B�`l�+z�]|���x��m�\�-[�����tw���j/^��=n!����wܼq���.�i���X!�ܘ���J�F�Z�|�<}Wzi}e	��!�\���;����暀����ɘ����in�������Zi~+����
aW�k��wwuNb�r�,[���%SA5��q	7�,�iz   �"�mM��vV�Z�_��?`J���;��	#s����/`^��ʀ�E�W�$�ilpr�H����������΢U�S��BG�6�̴$Q�T���*����8�D����~��u��sPP�K�[��iw=��RDQ%�aE���~6��K׀�Օ�v�鍹�v��mB<M������wژ+WI�����%=MG�1k��А`�[صf��/Rs����PZr⤁T�do�>E䆵�#����B��!��-���>ͺ�Y��"Y��@L̖�9�P��ب�ئ���0�W�ţ�6�d�]@���Z����-��&�-i-�b1��UJ4j�P�N����+�\�<��/�Ȍh)N�    IEND�B`�  l�PNG

   IHDR           szz�  3IDATx���OTg��`Z\b�E*Rh�Pl"�%@p�q�f�e�¾��@ղ�� ��!���XTA���T�ɴi�ml�<����51�/��7��y�y��g͚�U����3�X�������^i��<~��~yʽ�y��3!�222<EO^\ZZ���ĳ_����?x����=���؇� �jk�{�6�̓\��Ǣ^�\�Q\�y�h�+*+}�\��y����$7'�1�͘n�1s��%Tj�x]�/��sP�r||�3�����=�=���b2�0<<DKk�x ri4�]����p�|7���T������5.	�_77��{�nB����OWw�
TUU%F��C�xl��:��])�����}����<��������gq�P)2����t$���G��I�(�&א)@Qa:�m�T*9YY$%(hi�����bF�h�v��*�K�$D��b�6P\�CW[#��|b�d��H��V ,UFFF�P����Q��ɷ�-xyy-���7l�-""���ﹿ8Gxx8���A�RJ����"�F��I~|����9��Xb��$O���J����HPP�B�{3��Ls�3�swhl8���冔'�z   �G{kW��#CK��7c�&L��X\��zC-7F����N�]�899Qw�����N��Ya�/����g'�߱���)�$�=�W�ѣ���ͮ�}pp0Ey���g�T_Emuuߠq���t�֯�:׺:ɧnMQ��JIn^�%%�l�N�*�}*��V7��f�Z��|A��Z,������%�6��u"�C7�2tZ��8�{8r���J#�k�- ODC[[[B�{ �"��Z���Vi8^���뿢�c�7�Ş� ��G)�&m���-�p�pT..�QcӉ������ב���{�	�%6:��]�8\��BL�=PX2���(�$LD����#wlll��i 2�g����`�#�2t����ݷnu\vp��e��,1�B6���;����#��%7'S���"�J�>I(Iaa{���&)Q���s�+����T"�'Uvvv�����Y�mL��e�<6    IEND�B`�  j�PNG

   IHDR           szz�  1IDATx��iOTg��Ԗ,	5���e�4TLc�Q`�AE�� �:8(�̰8vFYG�a�m !����4�EAL���,��4�j���_ ��I���=9_��}���w�M���kb|��+,�/1��<*������g,>_`yi��Q��=7?Ttq������,o�~˛�oX{�&���U���ůD��������LM=dm�5���0vo���<C�#�ĳ�����Ƭc1=��Shkkc��8��tz�xUH�H����]&&&l���s��C�w��7n��Аq���nb����Bo_�n��`0������0�5F� 4xzH��Ԡ�^����BC�����gSr%[<�c)uf3:�%R�������H|BJE<��T� �gQ�U�
��=EJJ*r���'"Q�$�Rg��V<���T�����q2&E��FM��<��F����2����<�Bq�<N�	HM���Ŭ�]%3-�@�T&@x��s©�j52��B���\-�z   �zu)���^�;aTT��K,�2GDD����_�N߆��~<���<?�>,�W[%��>F��&�R�Lfx���O�y�������$�J)V)_�[��˗{
��=9y����Е�@_7U&{x01&��m��Z9���U`ii�,��.!�j͵H$J�t�47��"<9*���a�ފRZ>�c�:��p?����oA]}eF#&S��8��A*��*�@���J�:}��7Ӵe3��o���,]����'�l߱M�R0%e�Z�tv�����:����+�[����N�!ܺ�y�1��{��x9�q�%.ܶSi2`�6��Ձ��Ϫ�[	������p��đK۶Pj�S/İ����^������40��� b��8�k*�w��.#W� ��466^���Ɍ��'''¤���&��}!3�����0���b�'�s��f�wW"��p����|�ggg\]]�psuN���];���ό�����f�~�������|���yP��'=�11r��	�8JHh��-v3�Ҩ�#��㹱W���������c    IEND�B`�  ��PNG

   IHDR           szz�  HIDATx���O�wǽ�D�wA�	��9�	j̆�"TJ+�X
���Q�Z���ݰh@@���$�9ފ�0� �[\Щq�Ͳ��|�@�`�11�IN�\�����|�ϒ%oj���=�=ϟ>g��,�����V��k�ۮ�Lݟbn��c�<��6�����3>>�|�<���_��_��Fcc#�TUU1<<̕+�q��LOO311N[ۗ�k�`��C��yCqOoCCCtuv2:�=��8n�r��U�f�x]�h5�v}݅��bh�[����t:innfdd���~Z[���z8GK�P�ICC�0�::�QYYɵ�v���i���0��

�4�,*�[1[�X+�Ti-;L�q�x �cN�NRx� ���dj��%&�P(�P�b;z��L�x �!���z   �QVfD.�c0�'I����4�9A�<� ���P�T���LU
�JAA>E�z�&��{�i5�$F�$%9	ci1�Z-��l
�`�ͦ�l����o� b"#Q�����ޝ@z���\��ed������1�p?�'���,			���Pa.Ě"@*�r�f??�w��.Ϟ>^������@��~��쬧�}���>��\�t�K��v�������I$�N�1��s/fx����<�QM��t;��F�ZMrr2�D
�V�����df�kh@0�I��&��e�~�{�w�х������պ��]���4�r���<�q��8��s�u��wW066�g7�#C���=^T�U�V��8f�t� ��j�}N]�)�xg9���vw�������Khh��/b@@� <���1�R^�e�lo{P{҂������ گ���~�!��}P$Ɠ���e(wI��ɠ(v��o�t��GWZ/ �Ƌ�9
�@E�o	1$+��I%+sy˗R�WA�y���R����IاDE�"��"E�J)G�L��ϡI�xv\^� G��L&����v�V�|��!A�wG��#���o���"���P���_��-�ȤѤ)l�p[���/�������&8x��ylذ�����c���P����l�j1a*)$,<��;�,tc�$___�kq��]1��l۶� ��%�ǛJ��F}    IEND�B`�  ��PNG

   IHDR           szz�  fIDATx��]L�g�=�&n�%Kfb�&sʀM�M]�J�~���)�-C�?hH�Z��	
��
�����8�0⠀�T�N�L7��z��y�Ń%;فkM��9y��佯�~��{�I����]�E���qk�&���QS���2袧����nߺ͕�A��������?���������O�=��?���� ��={�#G���е!z����؀�̆e{�� R��-���t9�8q���n''N�����I}C=E�� t	���-�tvz   vr���n;�tt�x����::�����s _�mzv�mmm����jMM����k>J�p�QU�9 s��e˖1s�L�	z�۷a��Պ�؊�b����s �b��1���cT��i_�\�!QKI~6�Z�� ���l k��`H!"b��4��tj*K�NK�@���ul5e���HKO!#%��;��J�b��� �a�(�2̹[�)��z�d����ľ*zu~~~/{ 8  ���,��d��T�!�J���c?�\�*�l\�ۍT*�=��ڎB�@"	�t�	�4��6��*I��˥�����v�Z�(/�˦r��4n���=Ʈ���Μ>�,��������{��~Zf+�h�B����+�)N�ը����Zh&$$וK����?~�{w~���?
'$��N��hD�׮]��@�5��rpm�ŭ�c�\s�&�r��G�]t?ğ�V� v~�N���E7l�����7�sᜓ�K�1:���K�[�nح�b�1j����}�W����Tjs7��d�6����_����5{�낏���
�F�r2(�7RVj�d�v�2�=��h>�(��%mgN�.�3qUO�
��=�Ą8�Ց$'����2��7���J�ԗ����vN�j�U��=�f�"J)E�>��iD+��QN�B�X���N!g�\Z�#AAA����Z9c�/z�(Y��pT�b�)�X�M�t�(|}}�`���d�'��>��x!sߞ��<1��*���[Md���2`	�hV/�CЂ9�Z��i��ց��LFF*�P������wY�t���'J!!^�Y#C�R!Z�;h�q/���{�R)��J-Z��ٳ?����8�n�	u�    IEND�B`�  ÉPNG

   IHDR           szz�  �IDATx��L�u�ݲ�SˢaF�j���hY��"�s��8��~q��wp?9�;�D-Q�ɏ�d-�$�S��.��l�U$��b�����?�;�Z���gz   Ϟ����|����L��o]�=��N� }W�Q��S����_�p��� �ǭ�����A��^,V�7>/+�1z��ex��ёQ��c���Cnjjj�9@��΅�9r����n7׮�q���Xl��|&n0�ZZ[iw�sBX���.'�5�8�g8v�(y�y�sA��j=ъ�&A�Ч�hkk�^���������w 5�$7x���x��=ֈ�b���8��+�v�� +;��!!�:o�4=��B�ڱڬl-,��o�� �w �m��,߁)'mJ��T$R)R��\LE���4�� ��Š��0�J$@�Ƙ�(�b�:��R��C�ff ��9��q(���ofo��dy�T�� D�$'%b+ڊL.���h4`L�RQ^�^HKD����.�Y���8�8�����4���kQ�6/&E�A� 2Ұ��PVbf٢e3�Vd�cb��d�.�{�����?Q*�@<r��B�۫�)�M�M�?������ޏw�)D%�I1���=/+�V��b��ѣ�<��gMM��ř��n�UI	��1��\�L*![�����ss��;�an����~{���Fx'*j��^tt�[�'U<�����E�{�{g�����d��u��b0���U�+�#_7)z�]�f�	ι��@|7x��Y����}��%�Ȉ{�H��ם���P=��Oe��)�TWqxI��f\N]�N.�t�����h�n=�[��X�ī�����������(>��U�M���L��Fa��y��ߒ�g�Dhh(�Y�j�1`XD��r����0�|˔IO�L���:��ԌW ����/_�&�:5)���7�i�j%��M�T2��ɘ)�s�e�b����T̝;��K��D�(�4>e��7 �}�sO)�t1~~~�>�y�:fϞ͂���Hp�|�5���
�Z�b�ڔ�-��)lV)�X�����	^D�� ��Ŵ����n�a��{w9��x������6o{ʧ����9������C�z   �ӰV	�G�
w=鿱�3f�Ϛ�?g�+=����;���>&�     IEND�B`�  ʉPNG

   IHDR           szz�  �IDATx��mL�W���"�̐а��q3����0]1�P^kA(��Rii��A' FС(2���Y��+�`TT�Ȝ�)�̹�d�S�]�Oۇ�vf�Nrrs��y������gܸ��Y,-��+C~y�C���������\�z�����p�"='{���/u{p��T700����q����42JÞ=������sg9~��'{���yt���g8p� y���7�L�m�m���p��qN�Nb�����1�1��-���ܗ�^g���Sfe��
,��4448a:;;��:�����$��w��=�Ku�V0�-��}{5-��tt�S���} .dΜ9$J$��:�R)��SUUEA�*���u�(+� ����U�(i,�ˑ&%���@fz*����nXW\D�:�5&#qqq���"Nrb,�擗��>��eȃ_�h�G"I`� ��d�L����(�ձB��� mmm1��V�����6�W�eɗ#KMa��|H���fk�3� �o4�$>�������Aת������U���Ь�D�ӱ�` 5m9Y��=����jBB���ێt�T_�F�A���}{�� �Z����9::��@�Tʛ��"[�@q�����L��<��tZ*�6vg�<"""�
M&����c�pX���$¶T)�]_|*��o�1xT���	���/�7|��G��cc��!�
�s;��;Z�s}���b1�W.1|��;��t̻|s� �D�ȵK��w~��ӳ%22���/p����;�����s�}k�_�2����x���-}�!A��0;�������}4{O��i�o^�����~�� 2L{�ŵQQQ��]�l�јK���<�'=��@vl�f�b�: �z�D�a�k �ϟ/


�zk�+J)4�q�:��Sd2P^ZD�zk�1N�t��M%|z   l�E$Mxb�iӦ5��_��W��ΧE�V ���Jm:ٙ2�Q&��-�U)de� ��:|||��B�� -9����鯠�%��K�Ic��W���Z�I�IG�a�T?B���������!������m�-2���@&��ܲ(�C��\��3����/��f
��b��k������r�����}?�y3_b��Ag�ZG�p[�g�d��h��T��� �`�N���ƋD/v/��zj ����7���5$A�O    IEND�B`�  �PNG

   IHDR           szz�  �IDATx��L�e�]mj����@	Laci*HS��D �?<��〻�~� r`�z%������5�S��@祠��
PKg�By��?jk�vWk�={�}�Ϟ��y?������_֑&K��O6n�����h��r�3.}�MO�e�X�9w�«G�\��y���r��*���1��Ύ����:�� �yy�|n������h�� ��w�{�nR32\�<�dzf߾�X,Ξ=�ɓ���Zi;��Ν;���.��#��F��9�؈���e�����Tj�l6��b����ʪJ��GEQ�PO{{��'8d>D��&��Vq\�kj����#���|��ߡ�|3���h��UWc>l������ʌ������>]K�RIJj2ZĐ�F��a�[k?���r�:-��YȓdHerBBCH�"&"M�I|��tuu�jkk=�Ws�T�r�#:��D̫���ǊH\-�ݜtr�U��$?@E����TTT����V��Ő��@/�R��5�LEy�Q%)�z(�me%��@���h4R_[���9�,^�B.%w�u����h�r��D�Kֳt���;�cǪF�,%[��V�ak�_�2���>�f�������x��q̞5�7B��R���5ܻs��=�D$	;<Ѥ��,���bcc�s��S�����D"�E�Xj��/�/.z�%��>8�8�:W�z�7	��DDDi{��+�88����鉿z   �?�|}ab8� �[+�%0xo�����N�͘�4��i���B�r��wt]�����4�u��W����������MXXX���		�/��eg�ӭ�;z���w��?��jo7��o�0^�|y�Mh�ێ�I>v^9f5cF�G��=um2�t�Lk˧t�5s�^��#X�z��5l�PH��(5S [ͦ4�𬀒�)���a��#)^�E���������7�9df�Y��%M�z��F�S��L�
�(�R�RG�,�8'''�9���^HP�����'1���$�$1�m��Q(����� Q-�[E����������������ĉNL��²� �~�C
��*���D-<��5Q�
�Lqg�3�ލ)�n,X0���%�HS)�J
IS'Uo5yy���sΎ�Ns���ɓ��{���S�~��M�J		�̝�"η�����������K�,�w ��=�������    IEND�B`�  ��PNG

   IHDR           szz�  �IDATx��}L�uǭ���4kA!��u�b>5����ӝp�1�q��w���t�
� 5Q�BEQ��|���E�Ç��'�����mm�Q�����g����m��>�����~��a�u1�I8ą��}ϵ��9y�Wۯ0d v{�_�tw��}�>W:����4�";7��=tv��ȉ��i������6iD�gm{ill�H��C.^�������A]ݷ���Ha0�m6---r��~JKK������55[�Z�V: ]||���ijj���3�ڽˡF}�N�;*���ZS-���3��H��:��ʨ����_�g�jm%��T�)�`YN6���x{{���@jz*f�	��BE�JV,Mgͪ���u���b�@ͼ��J�Dz���,J��`sE9)>��|�6F���h,f=��I6�=��Ç}�kmul%a��S�ɠ'VK�5���јL\���R��Jѣ��z   N��ʒ���T����	F��"oI*q"�`���4RL�I:4��O/�޺�ڝ���JcYV&��XN������ϒ��D���������ϛo�g�܏\�b���u����h��Y&�5���{����x}����C���F�!,TA��:���WU,4������"-��=P(ܸ��@?��OD�8���NT*�4�_����L�AAAܼ���_�00�������<y����u����w*�9j����c����-t޺ɏ헱߽C�K���q}{��G��BH�F@@ g�5s⠍֖f.��g��w�����{<|�ã�:B.��m�R�_pa݋����i�������G8~��P�7�	��v�����ח�6��tu>�+��(!��1�������Q�)=���#�肭���s'� >>��y,'`�Ō5�$�f��%MOV�"�f.�jN� 7���hr�&&Lx�y
�d2,&��	�bըF>���1$i#H��"!6�D1ƪ�2g��ƍ˖���������}<�sW77��^���U�M�*�Oi|�?��
&	E&N|�I�2!�ۼ%��)�}���f3�K
X�2�U�+.�hT�)�H�)�v�$B���b�!��E�|]��}��rfϑ�/�th."S��4�H���D�"\5w�nB����Pݶ4$��    IEND�B`�  ��PNG

   IHDR           szz�  nIDATx��L�u�m�̜4�fSD@)hS���h�m5�Gw"����p�'��$H����]���	t`��H�J*`�z���?��K������g{����<���0�i<B��G��y������s��S��{�*O`hp��[�f��=�����Ӌ��$>DֆlM���s������=jkk�t�=t� ��FZ[O�s�G���9w���_��>B��ă��i�2��X,���̖�-T����3TW�b[E�x Q*�Hݾ:�DG��SM�hh��ĉ�Be��])���z   o-��@�JKK)//c�����KE�V�*��*� [h@///,X�&FMښ4R�R��H��`Y�ɔ����GN��pe�AAHH��B��`]��:R<��Y�$��MFj�!����2T�&B�!1C��8�V<�5i�(ÕI���OH@��&-QK�.
c�eD�x �����:2:z\� @�&'��W"�=�xMM;w���a�N���|����d�eA�����ቝ�l�g���AvF��p���d��Ơ�i���r�h���=RYY�\�B���]�6#{$�����{�㗾vϮ���J�����7A�RR�Y�i�!������������6�c��\��B��Uﻸ�x�2D·>�,��$=�$� �ō�� �����>��T*�$��/�+��꠫���}��E���y����<~��� ����_� ˷��gO��D�13&o/:�Oq���t}��}=޹e�1|h8�-�@���DR2u
�^���f�099y�0g�[�N 찜!F������F777
���Lc���6�'o�Rr�VS��$>��U�xj�����c\���p������V�<^�!%IG�NE����i���hY��� 	��/�9e�����vwww�A̝;Ud��~o�	���\%%L�*LF�&�*�lc��o���l�~�5˖�3g2cƫ�����u'��92�֖��_aڴi���U˗�zU �ί��� d逭�,�����\4a�1�f|�-���1�؎��W���|QQBQQ��6	6͒%���4���|F22Ra�`���_��®X�������7�Ǝ�S��    IEND�B`�  ��PNG

   IHDR           szz�  [IDATx��kL�g�]u�$�a3��F"�1q�S!P��hq�ȭ �K�i-��܆�z�W.�d���A@�"�P�3:��X\�e��=6��>L^�����$��9�9��s��q��eٙ3�z   ���k���1�����bbl��"n������3�3<�����O;A�.�IQPX@{�%��Ǹ><�Ӹ7�����������q�����;ʈ���� ���o9O�Z-D��������79p���K���������~jjNQ}�Z: �NGSs�������+tvuRU]E__/�g��9)���e�vD�����|ZBm]������q𠝣�B� 
�
���b���dff`���l�$wg.{�w�k1r�t�t %{K�]����lLF����r�)�u��Ӓ1�u��fgay�m�蒶�q�F4	qS4��s2d�ҥH5���Mb��,Qv֬,�!�NA���DB��7� ���IH�gW^Z]2�q"{c*;�&��.�ֈb�LNN&22�迻��K�����fy6���酓����#��kS��F���=�J�s*�c���|������1꠯��Z�f�+�T[ͩS'��g��{
��)���=f����㣢�����}�
�����$66�5>kF�U�ٔ&zl�����#��fb�)�{� E%n������l6�S�:�W�JEPP�XB���e����E������2�͉�G	����L������c�=_㈇�]�A��+|}����=�gݺu�>/��m��$���<�U}Fy�~��t�O���4�����:�[�%ZxmV	����ڑNF�c�NX��n��Y��2�r��3�'hin�r�jO�}/X�d	��!���'��CR�i�nғ�]�R)&����/�7>xy�!-Z��f%��0���$Do"1N�6��C"�W������O� �#z{{�
<==��Rl Z �7�F�%�+VH����Pq�n�����>>��UQ(�
���u����R������D�l��B�-{�����������=h4j�I|��U�V�92Bz����C2z�z�F�7�6@����/�����d��s�8q    IEND�B`�  j�PNG

  z    IHDR           szz�  1IDATx���O�U��E�J��jlڐ^H�V�e��Z&d�2�Ё�a�vX:��S:PdiӔ(�e(�L7�aQ/Z5��7&�5<��_�?��97����~�l��_�	뭾���{f��{C��������C�WXZpp{�"^��+����?>��~�?�dٱ���F���!�j��u�Ƭ}��ϦX���U��fF�V�(���h����f�K��sv�v;w��aph���~d2�x.�j5[��uю��X��hoog||����tuu���$@�\Nǵ�����L٦����u��m�/����/ǵ��כ�������.�������ڳ����0T(D��������i�Qg���B�U�a����<� ����2=yyj2��D�EZj�z+�R���@_V���e��rQ�ˉ��$��q�r��Uc�(F�R���P��~*��|J�z
���h��(����8]�%�X�h qqq(�����������D�ir��\i>G``��I�T*env���h����|s�Gc0�hŏa�D����w��gan���r�\		�'?K����aa��������4'81-\�l""��gɿyb�$-..ޞ���b��.�edd4����X7c�
�p�3�g�:1BPPujœ9����M�r=�Hmni��� Z�L�]��Z�9>����}L߳1?�W\��S&e��0A~o?���"���*!f�TU���NSC-&�����\�Ԉi�3��7���I��O��F�������g�����N��BC�)��44������������y�b�q������"{�	Ŷ��9A��34�R/8��l�О��+�@N<�&�W�1$�ǒ�L#�Ӕ�Ta�;��������{_ݱ��@��!K�#Q�r�f
��Yw�B}��a�R);]\\
 B��J���D��q��g��{�(��^!~cٹ�uv��E� "O�gϞ=����>%�İo��z   9 ��d�6�ڽ}c�:M6�t�tbc������A��<IHHxIt /��3���@�1p(,��G�ߍq����%��X��    IEND�B`�  e�PNG

   IHDR           szz�  ,IDATx�Ֆ}LSg�k�N5f ���i���B�X%mJӮ4tBJhצ0ڴ��vt���Ć�1� -+�!Ө���\��Ȍ����vL��ǒ�%;��}s�����sϽ�P(��N}���W`u3�턿Fx��b��NQ�f-�̈́8�>�[&�{�ߥ�63u����_�������]:� �ccW>���q |||ss/�߹s���^n��"�����N�L���k�/@���-���&��Ȱ�����s��__ ��=���̠e@ݠr��}x0u��<��O1yogg0q�::P)���XLFk>=�r؝�:}��h�m��r��q�ilx3h n���P�d(ɧ�Q̓����2�[Z����f5������E���q�فn� pՇ�g{q�oqA�E�J�$,+�
Ċ<�:��#�*%���x��0aT+1�������
��<oA� �J��TZ�QfCc[��Zz�����8p�mp�QUĜ�e��M�2����n 45i�r����.$��Vq�mf�	y(�ξ��+��2�/�9�b1�P�`@�P�h2bO|<�D1�4`3���t�Vnߺ�i�"S]�B/�!���.�󠪫GFT��i	ʑ����zxx(m��gj�o�"���@��"���@z33���$Bhja)e�U*�E_���]�D����1O�Mڵ�܌�2�Ǔۯ���71Γ��L/疢�i�K�Ew�
�V=�n_
�P�����V�~��0)H���i��݀�����^������Mp��p5*P##t˦�C)Iy9�G����*�!� \NM��M��e|ĆR�f��QX���J�����j����ϣ�Qp[��c�I���eӣ��V碀��.z   ��AI!��>���td< jT�@�N�����9I	m���\�������:�3�xl(e�+x(� $^El��՝;c>		��}� �?���ĥ��[~.�J���Y��h3@&��U�F��|/Fٱc� k�ˢA�2���2N)�f.�zq~�\b���o֖�t¥�O����h�̀UU�":�y}�̙���*V�t�V����q�ZN
���}���{W��]�'*�/(+x���^35���0B�|��o\?['�YVʥ��2�l����1ai��l�A4�k����E�O��Nb�1=*)f&�ޝ��.�24���C��5���G�O�8
���.�W���=���ɦ��������|8\)#U���b4���X,8,��5F((w�eR�Z���-���žt/%y���޽/��D���o�7��o�7�f    IEND�B`�  c�PNG

   IHDR           szz�  *IDATx��[L�u�I�mo:�23���2�6`PHǸL�ri�r-��B��P
��0�ld�Lf"0l���P���t��h����_�|�?�O�>��9�s�����*���j��w���c��]��ǣ�-�����=Xgdd�������cuy���=�N����_���Svv~�ɯ����-���c��"���LO�`~�+?~��/y��9;�;LLLP[���k�ɗ��feu��lm��������0��� 1ϥ˗�15���`c� ����x *�ꍉ�!���������M�~��_���c�W��;�|����h�v3�F�;������o`���ݔć�On������܄Vo���Aw� �mm��:�w��\UI��U<��B�ˋ���Q�������@�V���F[L�� ���qZ�����Ց�����@}C��0V���iqwwG.�7�9�P���;-�Ft�&J�5��+)�h���Q�((/U����� _<<<��j�⹵�D]�I�B� �.z  0�B+rs�H��Q! ��2��8-�0����m�Ef2��g��#��D��h_N���amdb��{zz�b:+'""��"%����`N�e��&$( SC5c}x{{�=��07�p22��jc�HO;KTT��A����.��J��L���1,&���dff���"((� ? �<E^^^�$|��'ve�c>����q�e1H$o�{�����Tt8�2�:ACC=9�l2#�x�]���D"1"$?'��#��^,\"+#�����}������>G����#����_�񵙙١�[��r�
#cc©�HOO.�������ͳ�j%z��V������'�t:��Ԑ��FFj2��L��<*ԅ8ڬ�{R��/�ZM��T���\x����Q�*Of6�_�ƴO:��N���,����8�(((8�o�K	&>ԗ���ݽ),���X�U%����D�'&��.܂�]&%%bk�`28t��� �-Fd�DG�P��si��+����/-8x𠟷�׏'#����H���0:"X4Kn�ǫشnmgLp]    IEND�B`�x